library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity filter_table is
	port(
		clk:  in  std_logic;
		addr: in  std_logic_vector(14 downto 0);
		data: out signed(17 downto 0)
	);
end filter_table;

architecture arch of filter_table is
	signal addr_d:  std_logic_vector(14 downto 11);
	signal addrardaddr:   std_logic_vector(15 downto 0);
	signal doado_00:  std_logic_vector(31 downto 0);
	signal dopadop_00: std_logic_vector(3 downto 0);
	signal doado_01:  std_logic_vector(31 downto 0);
	signal dopadop_01: std_logic_vector(3 downto 0);
	signal doado_02:  std_logic_vector(31 downto 0);
	signal dopadop_02: std_logic_vector(3 downto 0);
	signal doado_03:  std_logic_vector(31 downto 0);
	signal dopadop_03: std_logic_vector(3 downto 0);
	signal doado_04:  std_logic_vector(31 downto 0);
	signal dopadop_04: std_logic_vector(3 downto 0);
	signal doado_05:  std_logic_vector(31 downto 0);
	signal dopadop_05: std_logic_vector(3 downto 0);
	signal doado_06:  std_logic_vector(31 downto 0);
	signal dopadop_06: std_logic_vector(3 downto 0);
	signal doado_07:  std_logic_vector(31 downto 0);
	signal dopadop_07: std_logic_vector(3 downto 0);
	signal doado_08:  std_logic_vector(31 downto 0);
	signal dopadop_08: std_logic_vector(3 downto 0);
	signal doado_09:  std_logic_vector(31 downto 0);
	signal dopadop_09: std_logic_vector(3 downto 0);
	signal doado_10:  std_logic_vector(31 downto 0);
	signal dopadop_10: std_logic_vector(3 downto 0);
	signal doado_11:  std_logic_vector(31 downto 0);
	signal dopadop_11: std_logic_vector(3 downto 0);
	signal doado_12:  std_logic_vector(31 downto 0);
	signal dopadop_12: std_logic_vector(3 downto 0);
	signal doado_13:  std_logic_vector(31 downto 0);
	signal dopadop_13: std_logic_vector(3 downto 0);
	signal doado_14:  std_logic_vector(31 downto 0);
	signal dopadop_14: std_logic_vector(3 downto 0);
	signal doado_15:  std_logic_vector(31 downto 0);
	signal dopadop_15: std_logic_vector(3 downto 0);
begin
	addrardaddr(15)<='1';
	addrardaddr(14 downto 4)<=addr(10 downto 0);
	addrardaddr(3 downto 0)<=b"0000";
	process(clk)
	begin
		if (rising_edge(clk)) then
			addr_d<=addr(14 downto 11);
		end if;
	end process;
	with addr_d select data(15 downto 0)<=
		signed(doado_00(15 downto 0)) when b"0000",
		signed(doado_01(15 downto 0)) when b"0001",
		signed(doado_02(15 downto 0)) when b"0010",
		signed(doado_03(15 downto 0)) when b"0011",
		signed(doado_04(15 downto 0)) when b"0100",
		signed(doado_05(15 downto 0)) when b"0101",
		signed(doado_06(15 downto 0)) when b"0110",
		signed(doado_07(15 downto 0)) when b"0111",
		signed(doado_08(15 downto 0)) when b"1000",
		signed(doado_09(15 downto 0)) when b"1001",
		signed(doado_10(15 downto 0)) when b"1010",
		signed(doado_11(15 downto 0)) when b"1011",
		signed(doado_12(15 downto 0)) when b"1100",
		signed(doado_13(15 downto 0)) when b"1101",
		signed(doado_14(15 downto 0)) when b"1110",
		signed(doado_15(15 downto 0)) when others;
	with addr_d select data(17 downto 16)<=
		signed(dopadop_00(1 downto 0)) when b"0000",
		signed(dopadop_01(1 downto 0)) when b"0001",
		signed(dopadop_02(1 downto 0)) when b"0010",
		signed(dopadop_03(1 downto 0)) when b"0011",
		signed(dopadop_04(1 downto 0)) when b"0100",
		signed(dopadop_05(1 downto 0)) when b"0101",
		signed(dopadop_06(1 downto 0)) when b"0110",
		signed(dopadop_07(1 downto 0)) when b"0111",
		signed(dopadop_08(1 downto 0)) when b"1000",
		signed(dopadop_09(1 downto 0)) when b"1001",
		signed(dopadop_10(1 downto 0)) when b"1010",
		signed(dopadop_11(1 downto 0)) when b"1011",
		signed(dopadop_12(1 downto 0)) when b"1100",
		signed(dopadop_13(1 downto 0)) when b"1101",
		signed(dopadop_14(1 downto 0)) when b"1110",
		signed(dopadop_15(1 downto 0)) when others;
	mem_00: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_01=>X"0000000000000000000000000000000000000000000000000000000FFFFFFFFF",
		INITP_02=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000",
		INITP_04=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_05=>X"0000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_06=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_08=>X"000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_09=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_0A=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000",
		INITP_0B=>X"000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0C=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_0D=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000",
		INITP_0E=>X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0F=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_00=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_01=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_02=>X"FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_03=>X"FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_04=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9",
		INIT_05=>X"FFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFA",
		INIT_06=>X"FFFDFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFB",
		INIT_07=>X"FFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFD",
		INIT_08=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFE",
		INIT_09=>X"00010001000100000000000000000000000000000000000000000000FFFFFFFF",
		INIT_0A=>X"0002000200020002000200020002000100010001000100010001000100010001",
		INIT_0B=>X"0003000300030003000300030003000300030003000300030002000200020002",
		INIT_0C=>X"0005000500050004000400040004000400040004000400040004000400040004",
		INIT_0D=>X"0006000600060006000600050005000500050005000500050005000500050005",
		INIT_0E=>X"0007000700070007000700060006000600060006000600060006000600060006",
		INIT_0F=>X"0008000700070007000700070007000700070007000700070007000700070007",
		INIT_10=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_11=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_12=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_13=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_14=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_15=>X"0007000700070007000700070007000700070007000700080008000800080008",
		INIT_16=>X"0006000600060006000600060006000600070007000700070007000700070007",
		INIT_17=>X"0005000500050005000500050005000500050006000600060006000600060006",
		INIT_18=>X"0003000400040004000400040004000400040004000400040005000500050005",
		INIT_19=>X"0002000200020002000200020003000300030003000300030003000300030003",
		INIT_1A=>X"0000000000000001000100010001000100010001000100010002000200020002",
		INIT_1B=>X"FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000",
		INIT_1C=>X"FFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFE",
		INIT_1D=>X"FFFBFFFBFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFD",
		INIT_1E=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFB",
		INIT_1F=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_20=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_21=>X"FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_22=>X"FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5",
		INIT_23=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4",
		INIT_24=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3",
		INIT_25=>X"FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3",
		INIT_26=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF2FFF2",
		INIT_27=>X"FFF4FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3",
		INIT_28=>X"FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4",
		INIT_29=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5",
		INIT_2A=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF6FFF6",
		INIT_2B=>X"FFFBFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8",
		INIT_2C=>X"FFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFB",
		INIT_2D=>X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFE",
		INIT_2E=>X"0004000400030003000300030003000200020002000200010001000100010001",
		INIT_2F=>X"0007000700070007000700060006000600060005000500050005000400040004",
		INIT_30=>X"000B000B000B000B000A000A000A000A00090009000900090008000800080008",
		INIT_31=>X"000F000F000F000F000E000E000E000E000D000D000D000D000C000C000C000C",
		INIT_32=>X"0014001300130013001300120012001200120011001100110010001000100010",
		INIT_33=>X"0018001800170017001700160016001600160015001500150015001400140014",
		INIT_34=>X"001C001C001B001B001B001B001A001A001A001A001900190019001900180018",
		INIT_35=>X"002000200020001F001F001F001F001E001E001E001E001D001D001D001C001C",
		INIT_36=>X"0024002400240023002300230023002200220022002200210021002100210020",
		INIT_37=>X"0028002700270027002700270026002600260026002500250025002500240024",
		INIT_38=>X"002B002B002B002B002A002A002A002A00290029002900290029002800280028",
		INIT_39=>X"002E002E002E002E002E002D002D002D002D002D002C002C002C002C002C002B",
		INIT_3A=>X"0031003100310031003000300030003000300030002F002F002F002F002F002E",
		INIT_3B=>X"0033003300330033003300330032003200320032003200320032003100310031",
		INIT_3C=>X"0035003500350035003500350034003400340034003400340034003400340033",
		INIT_3D=>X"0036003600360036003600360036003600360036003600360035003500350035",
		INIT_3E=>X"0037003700370037003700370037003700370037003700370037003700370036",
		INIT_3F=>X"0038003700370037003700370037003700370037003700370037003700370037",
		INIT_40=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_41=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_42=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_43=>X"FFFCFFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFA",
		INIT_44=>X"FFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFC",
		INIT_45=>X"000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFE",
		INIT_46=>X"0002000200020002000200010001000100010001000100010000000000000000",
		INIT_47=>X"0004000400040004000400030003000300030003000300030003000200020002",
		INIT_48=>X"0006000600060005000500050005000500050005000500050004000400040004",
		INIT_49=>X"0007000700070007000700070007000600060006000600060006000600060006",
		INIT_4A=>X"0008000800080008000800080007000700070007000700070007000700070007",
		INIT_4B=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_4C=>X"0007000700070007000800080008000800080008000800080008000800080008",
		INIT_4D=>X"0006000600060007000700070007000700070007000700070007000700070007",
		INIT_4E=>X"0005000500050005000500050005000600060006000600060006000600060006",
		INIT_4F=>X"0003000300030003000300030004000400040004000400040004000400050005",
		INIT_50=>X"0001000100010001000100010001000200020002000200020002000200030003",
		INIT_51=>X"FFFEFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000",
		INIT_52=>X"FFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFE",
		INIT_53=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFCFFFC",
		INIT_54=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFFAFFFA",
		INIT_55=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_56=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_57=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_58=>X"FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_59=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_5A=>X"FFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_5B=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFA",
		INIT_5C=>X"FFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFD",
		INIT_5D=>X"000200020002000200010001000100010001000000000000000000000000FFFF",
		INIT_5E=>X"0005000500050004000400040004000400040003000300030003000300020002",
		INIT_5F=>X"0008000700070007000700070007000600060006000600060006000500050005",
		INIT_60=>X"000A000900090009000900090009000900090008000800080008000800080008",
		INIT_61=>X"000B000B000B000B000B000B000B000B000A000A000A000A000A000A000A000A",
		INIT_62=>X"000C000C000C000C000C000C000C000C000C000B000B000B000B000B000B000B",
		INIT_63=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C",
		INIT_64=>X"000A000B000B000B000B000B000B000B000B000B000B000B000B000B000B000C",
		INIT_65=>X"00090009000900090009000900090009000A000A000A000A000A000A000A000A",
		INIT_66=>X"0006000600060006000700070007000700070007000800080008000800080008",
		INIT_67=>X"0002000300030003000300030004000400040004000500050005000500050006",
		INIT_68=>X"FFFEFFFFFFFFFFFFFFFF00000000000000000001000100010001000200020002",
		INIT_69=>X"FFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFEFFFEFFFE",
		INIT_6A=>X"FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFA",
		INIT_6B=>X"FFF2FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6",
		INIT_6C=>X"FFEFFFEFFFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2",
		INIT_6D=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEF",
		INIT_6E=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFED",
		INIT_6F=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_70=>X"FFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFECFFECFFECFFEC",
		INIT_71=>X"FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEEFFEEFFEE",
		INIT_72=>X"FFF6FFF6FFF6FFF5FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF2FFF2FFF2FFF2",
		INIT_73=>X"FFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF7FFF7FFF7",
		INIT_74=>X"00050004000400030003000200020001000100000000FFFFFFFFFFFEFFFEFFFD",
		INIT_75=>X"000E000D000C000C000B000B000A000A00090008000800070007000600060005",
		INIT_76=>X"0017001700160015001500140014001300120012001100110010000F000F000E",
		INIT_77=>X"0022002100200020001F001E001E001D001C001C001B001B001A001900190018",
		INIT_78=>X"002C002B002B002A002900290028002700270026002500250024002400230022",
		INIT_79=>X"00360035003500340034003300320032003100300030002F002E002E002D002D",
		INIT_7A=>X"003F003F003E003E003D003C003C003B003B003A003A00390038003800370037",
		INIT_7B=>X"0047004700470046004600450045004400440043004200420041004100400040",
		INIT_7C=>X"004E004E004E004D004D004C004C004B004B004B004A004A0049004900480048",
		INIT_7D=>X"0053005300530053005200520052005100510051005000500050004F004F004F",
		INIT_7E=>X"0056005600560056005600560056005500550055005500550054005400540054",
		INIT_7F=>X"0058005700570057005700570057005700570057005700570057005700570057",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_00,
		DOPADOP=>dopadop_00,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_01: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_01=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000",
		INITP_03=>X"000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_04=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000",
		INITP_06=>X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_08=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000",
		INITP_09=>X"00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0A=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000",
		INITP_0B=>X"0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFF",
		INITP_0C=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000",
		INITP_0D=>X"00000000000000000000000000000000000000000000000000000FFFFFFFFFFF",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000",
		INITP_0F=>X"0000000000000000000000000000000000000000000000000000000000003FFF",
		INIT_00=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_01=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_02=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_03=>X"FFFCFFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFA",
		INIT_04=>X"FFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFC",
		INIT_05=>X"000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFE",
		INIT_06=>X"0002000200020002000200010001000100010001000100010000000000000000",
		INIT_07=>X"0004000400040004000400030003000300030003000300030003000200020002",
		INIT_08=>X"0006000600060005000500050005000500050005000500050004000400040004",
		INIT_09=>X"0007000700070007000700070007000600060006000600060006000600060006",
		INIT_0A=>X"0008000800080008000800080007000700070007000700070007000700070007",
		INIT_0B=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_0C=>X"0007000700070007000800080008000800080008000800080008000800080008",
		INIT_0D=>X"0006000600060007000700070007000700070007000700070007000700070007",
		INIT_0E=>X"0005000500050005000500050005000600060006000600060006000600060006",
		INIT_0F=>X"0003000300030003000300030004000400040004000400040004000400050005",
		INIT_10=>X"0001000100010001000100010001000200020002000200020002000200030003",
		INIT_11=>X"FFFEFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000",
		INIT_12=>X"FFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFE",
		INIT_13=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFCFFFC",
		INIT_14=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFFAFFFA",
		INIT_15=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_16=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_17=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_18=>X"FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_19=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_1A=>X"FFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_1B=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFA",
		INIT_1C=>X"FFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFD",
		INIT_1D=>X"000200020002000200010001000100010001000000000000000000000000FFFF",
		INIT_1E=>X"0005000500050004000400040004000400040003000300030003000300020002",
		INIT_1F=>X"0008000700070007000700070007000600060006000600060006000500050005",
		INIT_20=>X"000A000900090009000900090009000900090008000800080008000800080008",
		INIT_21=>X"000B000B000B000B000B000B000B000B000A000A000A000A000A000A000A000A",
		INIT_22=>X"000C000C000C000C000C000C000C000C000C000B000B000B000B000B000B000B",
		INIT_23=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C",
		INIT_24=>X"000A000B000B000B000B000B000B000B000B000B000B000B000B000B000B000C",
		INIT_25=>X"00090009000900090009000900090009000A000A000A000A000A000A000A000A",
		INIT_26=>X"0006000600060006000700070007000700070007000800080008000800080008",
		INIT_27=>X"0002000300030003000300030004000400040004000500050005000500050006",
		INIT_28=>X"FFFEFFFFFFFFFFFFFFFF00000000000000000001000100010001000200020002",
		INIT_29=>X"FFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFEFFFEFFFE",
		INIT_2A=>X"FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFA",
		INIT_2B=>X"FFF2FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6",
		INIT_2C=>X"FFEFFFEFFFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2",
		INIT_2D=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEF",
		INIT_2E=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFED",
		INIT_2F=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_30=>X"FFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFECFFECFFECFFEC",
		INIT_31=>X"FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEEFFEEFFEE",
		INIT_32=>X"FFF6FFF6FFF6FFF5FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF2FFF2FFF2FFF2",
		INIT_33=>X"FFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF7FFF7FFF7",
		INIT_34=>X"00050004000400030003000200020001000100000000FFFFFFFFFFFEFFFEFFFD",
		INIT_35=>X"000E000D000C000C000B000B000A000A00090008000800070007000600060005",
		INIT_36=>X"0017001700160015001500140014001300120012001100110010000F000F000E",
		INIT_37=>X"0022002100200020001F001E001E001D001C001C001B001B001A001900190018",
		INIT_38=>X"002C002B002B002A002900290028002700270026002500250024002400230022",
		INIT_39=>X"00360035003500340034003300320032003100300030002F002E002E002D002D",
		INIT_3A=>X"003F003F003E003E003D003C003C003B003B003A003A00390038003800370037",
		INIT_3B=>X"0047004700470046004600450045004400440043004200420041004100400040",
		INIT_3C=>X"004E004E004E004D004D004C004C004B004B004B004A004A0049004900480048",
		INIT_3D=>X"0053005300530053005200520052005100510051005000500050004F004F004F",
		INIT_3E=>X"0056005600560056005600560056005500550055005500550054005400540054",
		INIT_3F=>X"0058005700570057005700570057005700570057005700570057005700570057",
		INIT_40=>X"0007000700070007000700070007000700070007000700070007000700070007",
		INIT_41=>X"0005000500050005000500060006000600060006000600060006000700070007",
		INIT_42=>X"0002000200020003000300030003000300040004000400040004000400050005",
		INIT_43=>X"FFFFFFFFFFFFFFFF000000000000000000000001000100010001000100020002",
		INIT_44=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFF",
		INIT_45=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFB",
		INIT_46=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9",
		INIT_47=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8",
		INIT_48=>X"FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_49=>X"FFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9",
		INIT_4A=>X"FFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFB",
		INIT_4B=>X"000200020002000100010001000100000000000000000000FFFFFFFFFFFFFFFF",
		INIT_4C=>X"0005000500050004000400040004000400040003000300030003000300020002",
		INIT_4D=>X"0007000700070007000700070006000600060006000600060006000500050005",
		INIT_4E=>X"0008000800080008000800080008000800080008000800080008000700070007",
		INIT_4F=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_50=>X"0006000600060006000600060006000700070007000700070007000700070007",
		INIT_51=>X"0002000300030003000300040004000400040004000400050005000500050005",
		INIT_52=>X"FFFFFFFFFFFF0000000000000000000000010001000100010002000200020002",
		INIT_53=>X"FFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFF",
		INIT_54=>X"FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFB",
		INIT_55=>X"FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_56=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_57=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_58=>X"FFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_59=>X"FFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFA",
		INIT_5A=>X"00020002000200010001000100010000000000000000FFFFFFFFFFFFFFFFFFFE",
		INIT_5B=>X"0006000600060005000500050005000400040004000400030003000300030002",
		INIT_5C=>X"0009000900090009000800080008000800080007000700070007000700060006",
		INIT_5D=>X"000A000A000A000A000A000A000A000A000A000A000A000A0009000900090009",
		INIT_5E=>X"000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A",
		INIT_5F=>X"0008000800080008000800080009000900090009000900090009000A000A000A",
		INIT_60=>X"0004000400040004000500050005000600060006000600060007000700070007",
		INIT_61=>X"FFFFFFFF00000000000000000001000100010002000200020003000300030003",
		INIT_62=>X"FFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFEFFFF",
		INIT_63=>X"FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFA",
		INIT_64=>X"FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF5FFF6",
		INIT_65=>X"FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3",
		INIT_66=>X"FFF4FFF4FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF2",
		INIT_67=>X"FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF4FFF4FFF4",
		INIT_68=>X"FFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_69=>X"0003000300020002000200010001000000000000FFFFFFFFFFFEFFFEFFFEFFFD",
		INIT_6A=>X"0009000900090008000800080007000700060006000600050005000400040004",
		INIT_6B=>X"000E000E000E000E000D000D000D000D000C000C000C000B000B000B000A000A",
		INIT_6C=>X"001100110011001100110011001100100010001000100010000F000F000F000F",
		INIT_6D=>X"0011001100110011001100110012001200120012001200120012001100110011",
		INIT_6E=>X"000E000E000E000F000F000F000F001000100010001000100011001100110011",
		INIT_6F=>X"00080008000800090009000A000A000B000B000B000C000C000C000D000D000D",
		INIT_70=>X"FFFF000000000001000100020002000300030004000500050006000600070007",
		INIT_71=>X"FFF5FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFBFFFCFFFDFFFDFFFEFFFE",
		INIT_72=>X"FFECFFEDFFEDFFEEFFEEFFEFFFEFFFF0FFF1FFF1FFF2FFF2FFF3FFF4FFF4FFF5",
		INIT_73=>X"FFE5FFE5FFE6FFE6FFE7FFE7FFE7FFE8FFE8FFE9FFE9FFEAFFEAFFEBFFEBFFEC",
		INIT_74=>X"FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE3FFE3FFE3FFE3FFE4FFE4FFE4FFE4FFE5",
		INIT_75=>X"FFE3FFE3FFE3FFE3FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2",
		INIT_76=>X"FFEAFFEAFFE9FFE9FFE8FFE8FFE7FFE7FFE6FFE6FFE5FFE5FFE5FFE4FFE4FFE4",
		INIT_77=>X"FFF7FFF7FFF6FFF5FFF4FFF3FFF2FFF1FFF0FFEFFFEFFFEEFFEDFFECFFECFFEB",
		INIT_78=>X"000A00080007000600050004000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF8",
		INIT_79=>X"0020001F001D001C001A0019001700160014001300120010000F000E000C000B",
		INIT_7A=>X"003800370035003400320031002F002E002C002B002900270026002400230021",
		INIT_7B=>X"0051004F004E004C004B0049004800460045004300420040003F003D003B003A",
		INIT_7C=>X"006700650064006300620060005F005E005C005B005900580057005500540052",
		INIT_7D=>X"007800770076007500740073007200710070006F006E006D006C006A00690068",
		INIT_7E=>X"00840083008300820081008100800080007F007E007D007D007C007B007A0079",
		INIT_7F=>X"0088008700870087008700870087008700870086008600860085008500850084",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_01,
		DOPADOP=>dopadop_01,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_02: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000",
		INITP_01=>X"00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_02=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000",
		INITP_03=>X"0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFF",
		INITP_04=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000",
		INITP_05=>X"00000000000000000000000000000000000000000000000000000FFFFFFFFFFF",
		INITP_06=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000003FFF",
		INITP_08=>X"000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000",
		INITP_09=>X"FFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000",
		INITP_0A=>X"FFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
		INITP_0B=>X"0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0C=>X"0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000",
		INITP_0D=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFF",
		INITP_0F=>X"00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF",
		INIT_00=>X"0007000700070007000700070007000700070007000700070007000700070007",
		INIT_01=>X"0005000500050005000500060006000600060006000600060006000700070007",
		INIT_02=>X"0002000200020003000300030003000300040004000400040004000400050005",
		INIT_03=>X"FFFFFFFFFFFFFFFF000000000000000000000001000100010001000100020002",
		INIT_04=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFF",
		INIT_05=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFB",
		INIT_06=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9",
		INIT_07=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8",
		INIT_08=>X"FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_09=>X"FFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9",
		INIT_0A=>X"FFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFB",
		INIT_0B=>X"000200020002000100010001000100000000000000000000FFFFFFFFFFFFFFFF",
		INIT_0C=>X"0005000500050004000400040004000400040003000300030003000300020002",
		INIT_0D=>X"0007000700070007000700070006000600060006000600060006000500050005",
		INIT_0E=>X"0008000800080008000800080008000800080008000800080008000700070007",
		INIT_0F=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_10=>X"0006000600060006000600060006000700070007000700070007000700070007",
		INIT_11=>X"0002000300030003000300040004000400040004000400050005000500050005",
		INIT_12=>X"FFFFFFFFFFFF0000000000000000000000010001000100010002000200020002",
		INIT_13=>X"FFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFF",
		INIT_14=>X"FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFB",
		INIT_15=>X"FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_16=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_17=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_18=>X"FFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_19=>X"FFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFA",
		INIT_1A=>X"00020002000200010001000100010000000000000000FFFFFFFFFFFFFFFFFFFE",
		INIT_1B=>X"0006000600060005000500050005000400040004000400030003000300030002",
		INIT_1C=>X"0009000900090009000800080008000800080007000700070007000700060006",
		INIT_1D=>X"000A000A000A000A000A000A000A000A000A000A000A000A0009000900090009",
		INIT_1E=>X"000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A",
		INIT_1F=>X"0008000800080008000800080009000900090009000900090009000A000A000A",
		INIT_20=>X"0004000400040004000500050005000600060006000600060007000700070007",
		INIT_21=>X"FFFFFFFF00000000000000000001000100010002000200020003000300030003",
		INIT_22=>X"FFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFEFFFF",
		INIT_23=>X"FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFA",
		INIT_24=>X"FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF5FFF6",
		INIT_25=>X"FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3",
		INIT_26=>X"FFF4FFF4FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF2",
		INIT_27=>X"FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF4FFF4FFF4",
		INIT_28=>X"FFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_29=>X"0003000300020002000200010001000000000000FFFFFFFFFFFEFFFEFFFEFFFD",
		INIT_2A=>X"0009000900090008000800080007000700060006000600050005000400040004",
		INIT_2B=>X"000E000E000E000E000D000D000D000D000C000C000C000B000B000B000A000A",
		INIT_2C=>X"001100110011001100110011001100100010001000100010000F000F000F000F",
		INIT_2D=>X"0011001100110011001100110012001200120012001200120012001100110011",
		INIT_2E=>X"000E000E000E000F000F000F000F001000100010001000100011001100110011",
		INIT_2F=>X"00080008000800090009000A000A000B000B000B000C000C000C000D000D000D",
		INIT_30=>X"FFFF000000000001000100020002000300030004000500050006000600070007",
		INIT_31=>X"FFF5FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFBFFFCFFFDFFFDFFFEFFFE",
		INIT_32=>X"FFECFFEDFFEDFFEEFFEEFFEFFFEFFFF0FFF1FFF1FFF2FFF2FFF3FFF4FFF4FFF5",
		INIT_33=>X"FFE5FFE5FFE6FFE6FFE7FFE7FFE7FFE8FFE8FFE9FFE9FFEAFFEAFFEBFFEBFFEC",
		INIT_34=>X"FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE3FFE3FFE3FFE3FFE4FFE4FFE4FFE4FFE5",
		INIT_35=>X"FFE3FFE3FFE3FFE3FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2",
		INIT_36=>X"FFEAFFEAFFE9FFE9FFE8FFE8FFE7FFE7FFE6FFE6FFE5FFE5FFE5FFE4FFE4FFE4",
		INIT_37=>X"FFF7FFF7FFF6FFF5FFF4FFF3FFF2FFF1FFF0FFEFFFEFFFEEFFEDFFECFFECFFEB",
		INIT_38=>X"000A00080007000600050004000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF8",
		INIT_39=>X"0020001F001D001C001A0019001700160014001300120010000F000E000C000B",
		INIT_3A=>X"003800370035003400320031002F002E002C002B002900270026002400230021",
		INIT_3B=>X"0051004F004E004C004B0049004800460045004300420040003F003D003B003A",
		INIT_3C=>X"006700650064006300620060005F005E005C005B005900580057005500540052",
		INIT_3D=>X"007800770076007500740073007200710070006F006E006D006C006A00690068",
		INIT_3E=>X"00840083008300820081008100800080007F007E007D007D007C007B007A0079",
		INIT_3F=>X"0088008700870087008700870087008700870086008600860085008500850084",
		INIT_40=>X"0006000600060007000700070007000700070007000700070007000700070007",
		INIT_41=>X"0002000200030003000300040004000400040005000500050005000500060006",
		INIT_42=>X"FFFDFFFEFFFEFFFEFFFFFFFFFFFFFFFF00000000000000010001000100020002",
		INIT_43=>X"FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFD",
		INIT_44=>X"FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9",
		INIT_45=>X"FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7",
		INIT_46=>X"FFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9",
		INIT_47=>X"000100010000000000000000FFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFC",
		INIT_48=>X"0005000500050005000400040004000400030003000300030002000200020001",
		INIT_49=>X"0008000800080007000700070007000700070007000700060006000600060006",
		INIT_4A=>X"0007000700070007000700070008000800080008000800080008000800080008",
		INIT_4B=>X"0003000400040004000500050005000500050006000600060006000600070007",
		INIT_4C=>X"FFFEFFFFFFFFFFFF000000000000000100010001000200020002000300030003",
		INIT_4D=>X"FFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFE",
		INIT_4E=>X"FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFA",
		INIT_4F=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_50=>X"FFFBFFFBFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_51=>X"00000000FFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFCFFFBFFFB",
		INIT_52=>X"0005000500040004000400040003000300030002000200020001000100010000",
		INIT_53=>X"0008000800080008000800070007000700070007000700060006000600060005",
		INIT_54=>X"0008000800080008000900090009000900090009000900090009000800080008",
		INIT_55=>X"0005000500060006000600060007000700070007000700080008000800080008",
		INIT_56=>X"0000000000000001000100020002000200030003000300040004000400040005",
		INIT_57=>X"FFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFEFFFEFFFEFFFFFFFFFFFF",
		INIT_58=>X"FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFA",
		INIT_59=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_5A=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6",
		INIT_5B=>X"FFFEFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9",
		INIT_5C=>X"00050004000400040003000300020002000200010001000000000000FFFFFFFF",
		INIT_5D=>X"0009000900090009000800080008000800070007000700060006000600050005",
		INIT_5E=>X"000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A0009",
		INIT_5F=>X"000800080008000800090009000900090009000A000A000A000A000A000A000A",
		INIT_60=>X"0001000200020003000300040004000400050005000600060006000700070007",
		INIT_61=>X"FFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFFFFFF0000000000010001",
		INIT_62=>X"FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFFAFFFA",
		INIT_63=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5",
		INIT_64=>X"FFF6FFF5FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3FFF3FFF3FFF3FFF3",
		INIT_65=>X"FFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF6FFF6",
		INIT_66=>X"0005000400030003000200020001000100000000FFFFFFFFFFFEFFFEFFFDFFFD",
		INIT_67=>X"000B000B000B000A000A000A0009000900080008000700070006000600060005",
		INIT_68=>X"000E000E000E000E000E000E000E000E000E000D000D000D000D000C000C000C",
		INIT_69=>X"000C000C000D000D000D000D000E000E000E000E000E000E000E000E000E000E",
		INIT_6A=>X"0005000500060006000700070008000800090009000A000A000B000B000B000C",
		INIT_6B=>X"FFFBFFFBFFFCFFFCFFFDFFFEFFFEFFFF00000000000100020002000300030004",
		INIT_6C=>X"FFF1FFF2FFF2FFF3FFF3FFF4FFF5FFF5FFF6FFF6FFF7FFF7FFF8FFF9FFF9FFFA",
		INIT_6D=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF1FFF1",
		INIT_6E=>X"FFEFFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFED",
		INIT_6F=>X"FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF3FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFEF",
		INIT_70=>X"000400040003000200010000FFFFFFFEFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF8",
		INIT_71=>X"001100100010000F000E000D000D000C000B000A000900090008000700060005",
		INIT_72=>X"0019001900180018001800170017001600160015001500140014001300120012",
		INIT_73=>X"00180018001800190019001900190019001A001A001A001A0019001900190019",
		INIT_74=>X"000D000E000F0010001100110012001300140014001500150016001700170017",
		INIT_75=>X"FFFBFFFCFFFDFFFE000000010002000300040006000700080009000A000B000C",
		INIT_76=>X"FFE6FFE8FFE9FFEAFFEBFFECFFEEFFEFFFF0FFF2FFF3FFF4FFF6FFF7FFF8FFF9",
		INIT_77=>X"FFD7FFD8FFD9FFD9FFDAFFDBFFDCFFDDFFDEFFDFFFE0FFE1FFE2FFE3FFE4FFE5",
		INIT_78=>X"FFD5FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD5FFD5FFD5FFD6FFD6FFD7",
		INIT_79=>X"FFE3FFE2FFE1FFDFFFDEFFDDFFDCFFDBFFDAFFD9FFD8FFD7FFD7FFD6FFD6FFD5",
		INIT_7A=>X"00040002FFFFFFFDFFFBFFF8FFF6FFF4FFF2FFF0FFEEFFECFFEAFFE8FFE7FFE5",
		INIT_7B=>X"00330030002D002A002700240020001D001A001800150012000F000C000A0007",
		INIT_7C=>X"006800650062005E005B005800540051004E004A004700440040003D003A0037",
		INIT_7D=>X"0099009600940091008E008B008800850082007F007C007900750072006F006C",
		INIT_7E=>X"00BB00BA00B800B600B400B300B100AF00AC00AA00A800A600A300A1009E009C",
		INIT_7F=>X"00C800C700C700C700C700C600C600C500C400C400C300C200C100BF00BE00BD",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_02,
		DOPADOP=>dopadop_02,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_03: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000",
		INITP_01=>X"FFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000",
		INITP_02=>X"FFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
		INITP_03=>X"0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_04=>X"0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000",
		INITP_05=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000",
		INITP_06=>X"FFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFF",
		INITP_07=>X"00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF",
		INITP_08=>X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000",
		INITP_09=>X"FFFC0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF00000",
		INITP_0A=>X"FFFFFFFFFFFFC000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0B=>X"FFFFFFFFFFFFFFFFFFFFF0000000000000000000000000003FFFFFFFFFFFFFFF",
		INITP_0C=>X"00FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000003FFFFFF",
		INITP_0D=>X"00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000",
		INITP_0E=>X"00000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000",
		INITP_0F=>X"0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000",
		INIT_00=>X"0006000600060007000700070007000700070007000700070007000700070007",
		INIT_01=>X"0002000200030003000300040004000400040005000500050005000500060006",
		INIT_02=>X"FFFDFFFEFFFEFFFEFFFFFFFFFFFFFFFF00000000000000010001000100020002",
		INIT_03=>X"FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFD",
		INIT_04=>X"FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9",
		INIT_05=>X"FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7",
		INIT_06=>X"FFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9",
		INIT_07=>X"000100010000000000000000FFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFC",
		INIT_08=>X"0005000500050005000400040004000400030003000300030002000200020001",
		INIT_09=>X"0008000800080007000700070007000700070007000700060006000600060006",
		INIT_0A=>X"0007000700070007000700070008000800080008000800080008000800080008",
		INIT_0B=>X"0003000400040004000500050005000500050006000600060006000600070007",
		INIT_0C=>X"FFFEFFFFFFFFFFFF000000000000000100010001000200020002000300030003",
		INIT_0D=>X"FFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFE",
		INIT_0E=>X"FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFA",
		INIT_0F=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_10=>X"FFFBFFFBFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_11=>X"00000000FFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFCFFFBFFFB",
		INIT_12=>X"0005000500040004000400040003000300030002000200020001000100010000",
		INIT_13=>X"0008000800080008000800070007000700070007000700060006000600060005",
		INIT_14=>X"0008000800080008000900090009000900090009000900090009000800080008",
		INIT_15=>X"0005000500060006000600060007000700070007000700080008000800080008",
		INIT_16=>X"0000000000000001000100020002000200030003000300040004000400040005",
		INIT_17=>X"FFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFEFFFEFFFEFFFFFFFFFFFF",
		INIT_18=>X"FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFA",
		INIT_19=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_1A=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6",
		INIT_1B=>X"FFFEFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9",
		INIT_1C=>X"00050004000400040003000300020002000200010001000000000000FFFFFFFF",
		INIT_1D=>X"0009000900090009000800080008000800070007000700060006000600050005",
		INIT_1E=>X"000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A0009",
		INIT_1F=>X"000800080008000800090009000900090009000A000A000A000A000A000A000A",
		INIT_20=>X"0001000200020003000300040004000400050005000600060006000700070007",
		INIT_21=>X"FFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFFFFFF0000000000010001",
		INIT_22=>X"FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFFAFFFA",
		INIT_23=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5",
		INIT_24=>X"FFF6FFF5FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3FFF3FFF3FFF3FFF3",
		INIT_25=>X"FFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF6FFF6",
		INIT_26=>X"0005000400030003000200020001000100000000FFFFFFFFFFFEFFFEFFFDFFFD",
		INIT_27=>X"000B000B000B000A000A000A0009000900080008000700070006000600060005",
		INIT_28=>X"000E000E000E000E000E000E000E000E000E000D000D000D000D000C000C000C",
		INIT_29=>X"000C000C000D000D000D000D000E000E000E000E000E000E000E000E000E000E",
		INIT_2A=>X"0005000500060006000700070008000800090009000A000A000B000B000B000C",
		INIT_2B=>X"FFFBFFFBFFFCFFFCFFFDFFFEFFFEFFFF00000000000100020002000300030004",
		INIT_2C=>X"FFF1FFF2FFF2FFF3FFF3FFF4FFF5FFF5FFF6FFF6FFF7FFF7FFF8FFF9FFF9FFFA",
		INIT_2D=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF1FFF1",
		INIT_2E=>X"FFEFFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFED",
		INIT_2F=>X"FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF3FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFEF",
		INIT_30=>X"000400040003000200010000FFFFFFFEFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF8",
		INIT_31=>X"001100100010000F000E000D000D000C000B000A000900090008000700060005",
		INIT_32=>X"0019001900180018001800170017001600160015001500140014001300120012",
		INIT_33=>X"00180018001800190019001900190019001A001A001A001A0019001900190019",
		INIT_34=>X"000D000E000F0010001100110012001300140014001500150016001700170017",
		INIT_35=>X"FFFBFFFCFFFDFFFE000000010002000300040006000700080009000A000B000C",
		INIT_36=>X"FFE6FFE8FFE9FFEAFFEBFFECFFEEFFEFFFF0FFF2FFF3FFF4FFF6FFF7FFF8FFF9",
		INIT_37=>X"FFD7FFD8FFD9FFD9FFDAFFDBFFDCFFDDFFDEFFDFFFE0FFE1FFE2FFE3FFE4FFE5",
		INIT_38=>X"FFD5FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD5FFD5FFD5FFD6FFD6FFD7",
		INIT_39=>X"FFE3FFE2FFE1FFDFFFDEFFDDFFDCFFDBFFDAFFD9FFD8FFD7FFD7FFD6FFD6FFD5",
		INIT_3A=>X"00040002FFFFFFFDFFFBFFF8FFF6FFF4FFF2FFF0FFEEFFECFFEAFFE8FFE7FFE5",
		INIT_3B=>X"00330030002D002A002700240020001D001A001800150012000F000C000A0007",
		INIT_3C=>X"006800650062005E005B005800540051004E004A004700440040003D003A0037",
		INIT_3D=>X"0099009600940091008E008B008800850082007F007C007900750072006F006C",
		INIT_3E=>X"00BB00BA00B800B600B400B300B100AF00AC00AA00A800A600A300A1009E009C",
		INIT_3F=>X"00C800C700C700C700C700C600C600C500C400C400C300C200C100BF00BE00BD",
		INIT_40=>X"0004000500050005000600060006000600070007000700070007000700070007",
		INIT_41=>X"FFFEFFFEFFFEFFFFFFFF00000000000100010002000200020003000300040004",
		INIT_42=>X"FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFDFFFD",
		INIT_43=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_44=>X"FFFEFFFEFFFDFFFDFFFCFFFCFFFCFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF9",
		INIT_45=>X"0005000500040004000300030003000200020001000100000000FFFFFFFFFFFF",
		INIT_46=>X"0008000800080008000800070007000700070007000700060006000600060005",
		INIT_47=>X"0004000400050005000500060006000600070007000700070007000700070008",
		INIT_48=>X"FFFDFFFDFFFEFFFEFFFFFFFF0000000000010001000200020002000300030004",
		INIT_49=>X"FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFC",
		INIT_4A=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8",
		INIT_4B=>X"FFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFCFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9",
		INIT_4C=>X"000600050005000500040004000300030002000200020001000100000000FFFF",
		INIT_4D=>X"0008000800080008000800080008000800080007000700070007000700060006",
		INIT_4E=>X"0004000400050005000500060006000600070007000700070007000800080008",
		INIT_4F=>X"FFFCFFFDFFFDFFFEFFFEFFFFFFFF000000000001000100010002000200030003",
		INIT_50=>X"FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFC",
		INIT_51=>X"FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_52=>X"FFFFFFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFF9FFF9FFF9",
		INIT_53=>X"0007000600060005000500050004000400030003000200020001000100000000",
		INIT_54=>X"0008000900090009000900090009000800080008000800080008000700070007",
		INIT_55=>X"0003000400040005000500060006000600070007000700080008000800080008",
		INIT_56=>X"FFFBFFFCFFFCFFFDFFFDFFFEFFFEFFFFFFFF0000000000010001000200030003",
		INIT_57=>X"FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFB",
		INIT_58=>X"FFF8FFF8FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_59=>X"0000FFFFFFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF8",
		INIT_5A=>X"0008000700070007000600060005000500040004000300030002000200010001",
		INIT_5B=>X"0009000A000A000A000A000A000A000A000A0009000900090009000900080008",
		INIT_5C=>X"0003000400040005000500060006000700070008000800080009000900090009",
		INIT_5D=>X"FFFAFFFAFFFBFFFCFFFCFFFDFFFDFFFEFFFFFFFF000000000001000200020003",
		INIT_5E=>X"FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF8FFF8FFF8FFF9FFF9",
		INIT_5F=>X"FFF8FFF7FFF7FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF4FFF4FFF4FFF4",
		INIT_60=>X"000100000000FFFFFFFEFFFEFFFDFFFCFFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8",
		INIT_61=>X"000A000900090008000800080007000600060005000500040004000300020002",
		INIT_62=>X"000B000B000B000B000C000C000C000C000C000B000B000B000B000B000A000A",
		INIT_63=>X"000300040004000500060006000700070008000800090009000A000A000A000B",
		INIT_64=>X"FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFDFFFEFFFF00000000000100020002",
		INIT_65=>X"FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF4FFF4FFF4FFF5FFF5FFF6FFF6FFF7FFF7",
		INIT_66=>X"FFF6FFF6FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2",
		INIT_67=>X"0002000100010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8FFF7",
		INIT_68=>X"000D000C000C000B000B000A000A000900080008000700060005000500040003",
		INIT_69=>X"000E000E000E000E000F000F000F000F000F000F000F000E000E000E000E000D",
		INIT_6A=>X"000300040005000600060007000800090009000A000B000B000C000C000D000D",
		INIT_6B=>X"FFF5FFF6FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFEFFFF000000010002",
		INIT_6C=>X"FFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF1FFF1FFF2FFF3FFF3FFF4",
		INIT_6D=>X"FFF4FFF4FFF3FFF2FFF1FFF1FFF0FFF0FFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEE",
		INIT_6E=>X"00050004000300010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5",
		INIT_6F=>X"001300120012001100100010000F000E000D000C000B000A0009000800070006",
		INIT_70=>X"0013001300140014001400150015001500150015001500150014001400140013",
		INIT_71=>X"000300040006000700080009000A000B000C000D000E000F0010001100120012",
		INIT_72=>X"FFEEFFEFFFF0FFF1FFF3FFF4FFF5FFF7FFF8FFF9FFFBFFFCFFFEFFFF00000002",
		INIT_73=>X"FFE4FFE4FFE4FFE4FFE5FFE5FFE6FFE6FFE7FFE7FFE8FFE9FFEAFFEBFFECFFED",
		INIT_74=>X"FFEFFFEEFFEDFFECFFEBFFEAFFE9FFE8FFE7FFE6FFE6FFE5FFE5FFE5FFE4FFE4",
		INIT_75=>X"000B000900070005000300010000FFFEFFFCFFFAFFF9FFF7FFF5FFF4FFF2FFF1",
		INIT_76=>X"002200210020001F001E001D001B001A001800170015001300120010000E000C",
		INIT_77=>X"0022002300230024002500250025002600260026002600250025002400240023",
		INIT_78=>X"000300060008000B000D000F00110013001600170019001B001C001E001F0021",
		INIT_79=>X"FFD7FFDAFFDCFFDFFFE2FFE4FFE7FFEAFFEDFFF0FFF2FFF5FFF8FFFBFFFE0000",
		INIT_7A=>X"FFBFFFBFFFC0FFC0FFC1FFC2FFC4FFC5FFC6FFC8FFCAFFCCFFCEFFD0FFD2FFD5",
		INIT_7B=>X"FFD9FFD6FFD3FFD0FFCDFFCBFFC8FFC6FFC5FFC3FFC2FFC1FFC0FFC0FFBFFFBF",
		INIT_7C=>X"002C0025001F00190012000D00070001FFFCFFF7FFF2FFEDFFE9FFE5FFE0FFDD",
		INIT_7D=>X"009E0096008F0088008100790072006B0063005C0055004E0047004000390032",
		INIT_7E=>X"010000FC00F700F100EC00E600E000DA00D400CE00C700C100BA00B300AC00A5",
		INIT_7F=>X"01280127012701260125012401220120011D011B011801150111010D01090105",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_03,
		DOPADOP=>dopadop_03,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_04: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000",
		INITP_01=>X"FFFC0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF00000",
		INITP_02=>X"FFFFFFFFFFFFC000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_03=>X"FFFFFFFFFFFFFFFFFFFFF0000000000000000000000000003FFFFFFFFFFFFFFF",
		INITP_04=>X"00FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000003FFFFFF",
		INITP_05=>X"00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000",
		INITP_06=>X"00000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000",
		INITP_07=>X"0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000",
		INITP_08=>X"00000000000000FFFFFFFFFFFFFFFFFFFF00000000000000000000FFFFFFFFFF",
		INITP_09=>X"FFFFFFFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFFFFFF000000",
		INITP_0A=>X"FC00000000000000000003FFFFFFFFFFFFFFFFFFFC00000000000000000003FF",
		INITP_0B=>X"000003FFFFFFFFFFFFFFFFFFFC00000000000000000003FFFFFFFFFFFFFFFFFF",
		INITP_0C=>X"FFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFFFFFF000000000000000",
		INITP_0D=>X"0000000000000FFFFFFFFFFFFFFFFFFFF00000000000000000000FFFFFFFFFFF",
		INITP_0E=>X"FFFFFFFFFFFFFFFFC00000000000000000003FFFFFFFFFFFFFFFFFFFC0000000",
		INITP_0F=>X"000000000000000000003FFFFFFFFFFFFFFFFFFFC00000000000000000003FFF",
		INIT_00=>X"0004000500050005000600060006000600070007000700070007000700070007",
		INIT_01=>X"FFFEFFFEFFFEFFFFFFFF00000000000100010002000200020003000300040004",
		INIT_02=>X"FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFDFFFD",
		INIT_03=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_04=>X"FFFEFFFEFFFDFFFDFFFCFFFCFFFCFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF9",
		INIT_05=>X"0005000500040004000300030003000200020001000100000000FFFFFFFFFFFF",
		INIT_06=>X"0008000800080008000800070007000700070007000700060006000600060005",
		INIT_07=>X"0004000400050005000500060006000600070007000700070007000700070008",
		INIT_08=>X"FFFDFFFDFFFEFFFEFFFFFFFF0000000000010001000200020002000300030004",
		INIT_09=>X"FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFC",
		INIT_0A=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8",
		INIT_0B=>X"FFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFCFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9",
		INIT_0C=>X"000600050005000500040004000300030002000200020001000100000000FFFF",
		INIT_0D=>X"0008000800080008000800080008000800080007000700070007000700060006",
		INIT_0E=>X"0004000400050005000500060006000600070007000700070007000800080008",
		INIT_0F=>X"FFFCFFFDFFFDFFFEFFFEFFFFFFFF000000000001000100010002000200030003",
		INIT_10=>X"FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFC",
		INIT_11=>X"FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_12=>X"FFFFFFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFF9FFF9FFF9",
		INIT_13=>X"0007000600060005000500050004000400030003000200020001000100000000",
		INIT_14=>X"0008000900090009000900090009000800080008000800080008000700070007",
		INIT_15=>X"0003000400040005000500060006000600070007000700080008000800080008",
		INIT_16=>X"FFFBFFFCFFFCFFFDFFFDFFFEFFFEFFFFFFFF0000000000010001000200030003",
		INIT_17=>X"FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFB",
		INIT_18=>X"FFF8FFF8FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_19=>X"0000FFFFFFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF8",
		INIT_1A=>X"0008000700070007000600060005000500040004000300030002000200010001",
		INIT_1B=>X"0009000A000A000A000A000A000A000A000A0009000900090009000900080008",
		INIT_1C=>X"0003000400040005000500060006000700070008000800080009000900090009",
		INIT_1D=>X"FFFAFFFAFFFBFFFCFFFCFFFDFFFDFFFEFFFFFFFF000000000001000200020003",
		INIT_1E=>X"FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF8FFF8FFF8FFF9FFF9",
		INIT_1F=>X"FFF8FFF7FFF7FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF4FFF4FFF4FFF4",
		INIT_20=>X"000100000000FFFFFFFEFFFEFFFDFFFCFFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8",
		INIT_21=>X"000A000900090008000800080007000600060005000500040004000300020002",
		INIT_22=>X"000B000B000B000B000C000C000C000C000C000B000B000B000B000B000A000A",
		INIT_23=>X"000300040004000500060006000700070008000800090009000A000A000A000B",
		INIT_24=>X"FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFDFFFEFFFF00000000000100020002",
		INIT_25=>X"FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF4FFF4FFF4FFF5FFF5FFF6FFF6FFF7FFF7",
		INIT_26=>X"FFF6FFF6FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2",
		INIT_27=>X"0002000100010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8FFF7",
		INIT_28=>X"000D000C000C000B000B000A000A000900080008000700060005000500040003",
		INIT_29=>X"000E000E000E000E000F000F000F000F000F000F000F000E000E000E000E000D",
		INIT_2A=>X"000300040005000600060007000800090009000A000B000B000C000C000D000D",
		INIT_2B=>X"FFF5FFF6FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFEFFFF000000010002",
		INIT_2C=>X"FFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF1FFF1FFF2FFF3FFF3FFF4",
		INIT_2D=>X"FFF4FFF4FFF3FFF2FFF1FFF1FFF0FFF0FFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEE",
		INIT_2E=>X"00050004000300010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5",
		INIT_2F=>X"001300120012001100100010000F000E000D000C000B000A0009000800070006",
		INIT_30=>X"0013001300140014001400150015001500150015001500150014001400140013",
		INIT_31=>X"000300040006000700080009000A000B000C000D000E000F0010001100120012",
		INIT_32=>X"FFEEFFEFFFF0FFF1FFF3FFF4FFF5FFF7FFF8FFF9FFFBFFFCFFFEFFFF00000002",
		INIT_33=>X"FFE4FFE4FFE4FFE4FFE5FFE5FFE6FFE6FFE7FFE7FFE8FFE9FFEAFFEBFFECFFED",
		INIT_34=>X"FFEFFFEEFFEDFFECFFEBFFEAFFE9FFE8FFE7FFE6FFE6FFE5FFE5FFE5FFE4FFE4",
		INIT_35=>X"000B000900070005000300010000FFFEFFFCFFFAFFF9FFF7FFF5FFF4FFF2FFF1",
		INIT_36=>X"002200210020001F001E001D001B001A001800170015001300120010000E000C",
		INIT_37=>X"0022002300230024002500250025002600260026002600250025002400240023",
		INIT_38=>X"000300060008000B000D000F00110013001600170019001B001C001E001F0021",
		INIT_39=>X"FFD7FFDAFFDCFFDFFFE2FFE4FFE7FFEAFFEDFFF0FFF2FFF5FFF8FFFBFFFE0000",
		INIT_3A=>X"FFBFFFBFFFC0FFC0FFC1FFC2FFC4FFC5FFC6FFC8FFCAFFCCFFCEFFD0FFD2FFD5",
		INIT_3B=>X"FFD9FFD6FFD3FFD0FFCDFFCBFFC8FFC6FFC5FFC3FFC2FFC1FFC0FFC0FFBFFFBF",
		INIT_3C=>X"002C0025001F00190012000D00070001FFFCFFF7FFF2FFEDFFE9FFE5FFE0FFDD",
		INIT_3D=>X"009E0096008F0088008100790072006B0063005C0055004E0047004000390032",
		INIT_3E=>X"010000FC00F700F100EC00E600E000DA00D400CE00C700C100BA00B300AC00A5",
		INIT_3F=>X"01280127012701260125012401220120011D011B011801150111010D01090105",
		INIT_40=>X"FFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_41=>X"000600060005000500040004000300030002000100010000FFFFFFFFFFFEFFFE",
		INIT_42=>X"0006000600070007000700070007000700080007000700070007000700070006",
		INIT_43=>X"FFFDFFFEFFFEFFFF000000000001000200020003000300040004000500050006",
		INIT_44=>X"FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFD",
		INIT_45=>X"FFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF7",
		INIT_46=>X"000600050005000500040004000300020002000100010000FFFFFFFFFFFEFFFD",
		INIT_47=>X"0006000700070007000700070008000800080008000700070007000700070006",
		INIT_48=>X"FFFDFFFEFFFFFFFF000000000001000200020003000400040005000500050006",
		INIT_49=>X"FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFAFFFBFFFCFFFCFFFD",
		INIT_4A=>X"FFFDFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF7FFF7FFF7",
		INIT_4B=>X"000600060005000500040003000300020002000100000000FFFFFFFEFFFEFFFD",
		INIT_4C=>X"0007000700070007000800080008000800080008000800080007000700070006",
		INIT_4D=>X"FFFDFFFEFFFFFFFF000000010001000200030003000400040005000500060006",
		INIT_4E=>X"FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFBFFFCFFFCFFFD",
		INIT_4F=>X"FFFCFFFCFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7",
		INIT_50=>X"00060006000500050004000300030002000200010000FFFFFFFFFFFEFFFDFFFD",
		INIT_51=>X"0007000700080008000800080008000800080008000800080008000700070007",
		INIT_52=>X"FFFEFFFEFFFF0000000000010002000200030004000400050005000600060007",
		INIT_53=>X"FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFCFFFCFFFD",
		INIT_54=>X"FFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF6FFF6FFF6",
		INIT_55=>X"00060006000500050004000300030002000100010000FFFFFFFFFFFEFFFDFFFC",
		INIT_56=>X"0008000800080009000900090009000900090009000900080008000800070007",
		INIT_57=>X"FFFEFFFEFFFF0000000100010002000300030004000500050006000600070007",
		INIT_58=>X"FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFBFFFCFFFD",
		INIT_59=>X"FFFBFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_5A=>X"00070006000600050004000400030002000100010000FFFFFFFEFFFDFFFDFFFC",
		INIT_5B=>X"0009000900090009000A000A000A000A000A000A000900090009000800080007",
		INIT_5C=>X"FFFEFFFFFFFF0000000100020003000300040005000500060007000700080008",
		INIT_5D=>X"FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFBFFFBFFFCFFFD",
		INIT_5E=>X"FFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF5",
		INIT_5F=>X"00080007000600050005000400030002000100000000FFFFFFFEFFFDFFFCFFFB",
		INIT_60=>X"000A000A000B000B000B000B000B000B000B000B000A000A000A000900090008",
		INIT_61=>X"FFFEFFFF00000001000100020003000400050006000600070008000800090009",
		INIT_62=>X"FFF3FFF4FFF4FFF4FFF5FFF5FFF6FFF6FFF7FFF8FFF9FFF9FFFAFFFBFFFCFFFD",
		INIT_63=>X"FFFAFFF9FFF8FFF7FFF6FFF6FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF3FFF3",
		INIT_64=>X"0008000800070006000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFA",
		INIT_65=>X"000C000C000C000D000D000D000D000D000C000C000C000B000B000A000A0009",
		INIT_66=>X"FFFEFFFF00000001000200030004000500060007000800090009000A000B000B",
		INIT_67=>X"FFF1FFF2FFF2FFF3FFF3FFF4FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFD",
		INIT_68=>X"FFF8FFF7FFF6FFF5FFF5FFF4FFF3FFF3FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF1",
		INIT_69=>X"000A000900080007000600050004000200010000FFFFFFFEFFFCFFFBFFFAFFF9",
		INIT_6A=>X"000E000F000F000F000F0010000F000F000F000F000E000E000D000C000C000B",
		INIT_6B=>X"FFFEFFFF00000002000300040006000700080009000A000B000C000D000D000E",
		INIT_6C=>X"FFEEFFEFFFEFFFF0FFF0FFF1FFF2FFF3FFF4FFF5FFF6FFF7FFF9FFFAFFFBFFFD",
		INIT_6D=>X"FFF6FFF5FFF4FFF3FFF2FFF1FFF0FFEFFFEFFFEEFFEEFFEEFFEEFFEEFFEEFFEE",
		INIT_6E=>X"000C000B000A0008000700060004000300010000FFFEFFFDFFFBFFFAFFF8FFF7",
		INIT_6F=>X"00130013001400140014001400140014001300130012001100110010000F000E",
		INIT_70=>X"FFFE0000000100030005000600080009000B000C000D000F0010001100110012",
		INIT_71=>X"FFE8FFE9FFEAFFEBFFECFFEDFFEEFFEFFFF1FFF2FFF4FFF5FFF7FFF9FFFAFFFC",
		INIT_72=>X"FFF2FFF0FFEFFFEDFFECFFEBFFEAFFE9FFE9FFE8FFE8FFE7FFE7FFE7FFE8FFE8",
		INIT_73=>X"0011000F000D000B00090007000500030001FFFFFFFDFFFBFFF9FFF7FFF5FFF4",
		INIT_74=>X"001B001C001D001D001D001D001C001C001B001A001A00180017001600140013",
		INIT_75=>X"FFFE0000000300050008000A000C000F001100130014001600170019001A001B",
		INIT_76=>X"FFDCFFDDFFDFFFE0FFE2FFE4FFE6FFE8FFEAFFECFFEFFFF1FFF4FFF6FFF9FFFB",
		INIT_77=>X"FFE9FFE6FFE4FFE2FFE0FFDFFFDDFFDCFFDBFFDBFFDAFFDAFFDAFFDAFFDBFFDB",
		INIT_78=>X"001C001900160012000F000C000800050001FFFEFFFAFFF7FFF4FFF1FFEEFFEB",
		INIT_79=>X"003300340034003400340033003200310030002E002C002A002800250022001F",
		INIT_7A=>X"FFFE00030008000D00110016001A001E002100240027002A002D002F00300032",
		INIT_7B=>X"FFB1FFB5FFB8FFBCFFC0FFC5FFCAFFCEFFD4FFD9FFDEFFE3FFE9FFEEFFF3FFF9",
		INIT_7C=>X"FFC1FFBCFFB7FFB3FFAFFFACFFAAFFA8FFA7FFA7FFA7FFA7FFA8FFAAFFACFFAF",
		INIT_7D=>X"006100530047003A002E00220017000C0001FFF7FFEEFFE5FFDCFFD5FFCDFFC7",
		INIT_7E=>X"01350129011D0111010400F700EA00DC00CF00C100B300A500970089007C006E",
		INIT_7F=>X"01980197019601940191018D01890183017D0177016F0167015E0155014B0140",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_04,
		DOPADOP=>dopadop_04,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_05: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"00000000000000FFFFFFFFFFFFFFFFFFFF00000000000000000000FFFFFFFFFF",
		INITP_01=>X"FFFFFFFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFFFFFF000000",
		INITP_02=>X"FC00000000000000000003FFFFFFFFFFFFFFFFFFFC00000000000000000003FF",
		INITP_03=>X"000003FFFFFFFFFFFFFFFFFFFC00000000000000000003FFFFFFFFFFFFFFFFFF",
		INITP_04=>X"FFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFFFFFF000000000000000",
		INITP_05=>X"0000000000000FFFFFFFFFFFFFFFFFFFF00000000000000000000FFFFFFFFFFF",
		INITP_06=>X"FFFFFFFFFFFFFFFFC00000000000000000003FFFFFFFFFFFFFFFFFFFC0000000",
		INITP_07=>X"000000000000000000003FFFFFFFFFFFFFFFFFFFC00000000000000000003FFF",
		INITP_08=>X"F00000000000000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF0000000",
		INITP_09=>X"FFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFF",
		INITP_0A=>X"000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000000FFFFF",
		INITP_0B=>X"00000000000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000",
		INITP_0C=>X"FFFFC00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC000",
		INITP_0D=>X"FFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFF",
		INITP_0E=>X"0000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC00000000000003F",
		INITP_0F=>X"000000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC0000000",
		INIT_00=>X"FFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_01=>X"000600060005000500040004000300030002000100010000FFFFFFFFFFFEFFFE",
		INIT_02=>X"0006000600070007000700070007000700080007000700070007000700070006",
		INIT_03=>X"FFFDFFFEFFFEFFFF000000000001000200020003000300040004000500050006",
		INIT_04=>X"FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFD",
		INIT_05=>X"FFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF7",
		INIT_06=>X"000600050005000500040004000300020002000100010000FFFFFFFFFFFEFFFD",
		INIT_07=>X"0006000700070007000700070008000800080008000700070007000700070006",
		INIT_08=>X"FFFDFFFEFFFFFFFF000000000001000200020003000400040005000500050006",
		INIT_09=>X"FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFAFFFBFFFCFFFCFFFD",
		INIT_0A=>X"FFFDFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF7FFF7FFF7",
		INIT_0B=>X"000600060005000500040003000300020002000100000000FFFFFFFEFFFEFFFD",
		INIT_0C=>X"0007000700070007000800080008000800080008000800080007000700070006",
		INIT_0D=>X"FFFDFFFEFFFFFFFF000000010001000200030003000400040005000500060006",
		INIT_0E=>X"FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFBFFFCFFFCFFFD",
		INIT_0F=>X"FFFCFFFCFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7",
		INIT_10=>X"00060006000500050004000300030002000200010000FFFFFFFFFFFEFFFDFFFD",
		INIT_11=>X"0007000700080008000800080008000800080008000800080008000700070007",
		INIT_12=>X"FFFEFFFEFFFF0000000000010002000200030004000400050005000600060007",
		INIT_13=>X"FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFCFFFCFFFD",
		INIT_14=>X"FFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF6FFF6FFF6",
		INIT_15=>X"00060006000500050004000300030002000100010000FFFFFFFFFFFEFFFDFFFC",
		INIT_16=>X"0008000800080009000900090009000900090009000900080008000800070007",
		INIT_17=>X"FFFEFFFEFFFF0000000100010002000300030004000500050006000600070007",
		INIT_18=>X"FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFBFFFCFFFD",
		INIT_19=>X"FFFBFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_1A=>X"00070006000600050004000400030002000100010000FFFFFFFEFFFDFFFDFFFC",
		INIT_1B=>X"0009000900090009000A000A000A000A000A000A000900090009000800080007",
		INIT_1C=>X"FFFEFFFFFFFF0000000100020003000300040005000500060007000700080008",
		INIT_1D=>X"FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFBFFFBFFFCFFFD",
		INIT_1E=>X"FFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF5",
		INIT_1F=>X"00080007000600050005000400030002000100000000FFFFFFFEFFFDFFFCFFFB",
		INIT_20=>X"000A000A000B000B000B000B000B000B000B000B000A000A000A000900090008",
		INIT_21=>X"FFFEFFFF00000001000100020003000400050006000600070008000800090009",
		INIT_22=>X"FFF3FFF4FFF4FFF4FFF5FFF5FFF6FFF6FFF7FFF8FFF9FFF9FFFAFFFBFFFCFFFD",
		INIT_23=>X"FFFAFFF9FFF8FFF7FFF6FFF6FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF3FFF3",
		INIT_24=>X"0008000800070006000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFA",
		INIT_25=>X"000C000C000C000D000D000D000D000D000C000C000C000B000B000A000A0009",
		INIT_26=>X"FFFEFFFF00000001000200030004000500060007000800090009000A000B000B",
		INIT_27=>X"FFF1FFF2FFF2FFF3FFF3FFF4FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFD",
		INIT_28=>X"FFF8FFF7FFF6FFF5FFF5FFF4FFF3FFF3FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF1",
		INIT_29=>X"000A000900080007000600050004000200010000FFFFFFFEFFFCFFFBFFFAFFF9",
		INIT_2A=>X"000E000F000F000F000F0010000F000F000F000F000E000E000D000C000C000B",
		INIT_2B=>X"FFFEFFFF00000002000300040006000700080009000A000B000C000D000D000E",
		INIT_2C=>X"FFEEFFEFFFEFFFF0FFF0FFF1FFF2FFF3FFF4FFF5FFF6FFF7FFF9FFFAFFFBFFFD",
		INIT_2D=>X"FFF6FFF5FFF4FFF3FFF2FFF1FFF0FFEFFFEFFFEEFFEEFFEEFFEEFFEEFFEEFFEE",
		INIT_2E=>X"000C000B000A0008000700060004000300010000FFFEFFFDFFFBFFFAFFF8FFF7",
		INIT_2F=>X"00130013001400140014001400140014001300130012001100110010000F000E",
		INIT_30=>X"FFFE0000000100030005000600080009000B000C000D000F0010001100110012",
		INIT_31=>X"FFE8FFE9FFEAFFEBFFECFFEDFFEEFFEFFFF1FFF2FFF4FFF5FFF7FFF9FFFAFFFC",
		INIT_32=>X"FFF2FFF0FFEFFFEDFFECFFEBFFEAFFE9FFE9FFE8FFE8FFE7FFE7FFE7FFE8FFE8",
		INIT_33=>X"0011000F000D000B00090007000500030001FFFFFFFDFFFBFFF9FFF7FFF5FFF4",
		INIT_34=>X"001B001C001D001D001D001D001C001C001B001A001A00180017001600140013",
		INIT_35=>X"FFFE0000000300050008000A000C000F001100130014001600170019001A001B",
		INIT_36=>X"FFDCFFDDFFDFFFE0FFE2FFE4FFE6FFE8FFEAFFECFFEFFFF1FFF4FFF6FFF9FFFB",
		INIT_37=>X"FFE9FFE6FFE4FFE2FFE0FFDFFFDDFFDCFFDBFFDBFFDAFFDAFFDAFFDAFFDBFFDB",
		INIT_38=>X"001C001900160012000F000C000800050001FFFEFFFAFFF7FFF4FFF1FFEEFFEB",
		INIT_39=>X"003300340034003400340033003200310030002E002C002A002800250022001F",
		INIT_3A=>X"FFFE00030008000D00110016001A001E002100240027002A002D002F00300032",
		INIT_3B=>X"FFB1FFB5FFB8FFBCFFC0FFC5FFCAFFCEFFD4FFD9FFDEFFE3FFE9FFEEFFF3FFF9",
		INIT_3C=>X"FFC1FFBCFFB7FFB3FFAFFFACFFAAFFA8FFA7FFA7FFA7FFA7FFA8FFAAFFACFFAF",
		INIT_3D=>X"006100530047003A002E00220017000C0001FFF7FFEEFFE5FFDCFFD5FFCDFFC7",
		INIT_3E=>X"01350129011D0111010400F700EA00DC00CF00C100B300A500970089007C006E",
		INIT_3F=>X"01980197019601940191018D01890183017D0177016F0167015E0155014B0140",
		INIT_40=>X"FFFEFFFF00000000000100020003000400040005000600060007000700070007",
		INIT_41=>X"FFF8FFF8FFF8FFF8FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFD",
		INIT_42=>X"000400040003000200010000FFFFFFFFFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF9",
		INIT_43=>X"0005000500060006000700070007000700080007000700070007000600060005",
		INIT_44=>X"FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFEFFFF000000010001000200030004",
		INIT_45=>X"FFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF9FFF8FFF8FFF8FFF7FFF7FFF8FFF8FFF8",
		INIT_46=>X"00080008000700070007000600060005000400040003000200010000FFFFFFFE",
		INIT_47=>X"FFFEFFFF00000001000200020003000400050005000600060007000700070008",
		INIT_48=>X"FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFD",
		INIT_49=>X"000400040003000200010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFFAFFF9FFF8",
		INIT_4A=>X"0005000600060007000700070008000800080008000700070007000600060005",
		INIT_4B=>X"FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFEFFFF000000010002000300030004",
		INIT_4C=>X"FFFDFFFCFFFCFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF8",
		INIT_4D=>X"00080008000800070007000600060005000400040003000200010000FFFFFFFE",
		INIT_4E=>X"FFFEFFFF00000001000200030004000400050006000600070007000800080008",
		INIT_4F=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFFAFFFBFFFBFFFCFFFD",
		INIT_50=>X"000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8",
		INIT_51=>X"0005000600070007000800080008000800080008000800080007000700060005",
		INIT_52=>X"FFF8FFF8FFF9FFFAFFFAFFFBFFFCFFFDFFFEFFFF000000010002000300040005",
		INIT_53=>X"FFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_54=>X"00090009000800080007000700060005000500040003000200010000FFFFFFFE",
		INIT_55=>X"FFFEFFFF00000001000200030004000500060007000700080008000800090009",
		INIT_56=>X"FFF7FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF9FFF9FFFAFFFBFFFCFFFD",
		INIT_57=>X"000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF7",
		INIT_58=>X"0006000700080008000900090009000900090009000900080008000700070006",
		INIT_59=>X"FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF000000010003000400050005",
		INIT_5A=>X"FFFCFFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF6FFF6FFF6FFF5FFF6FFF6FFF6FFF6",
		INIT_5B=>X"000A000A000900090008000800070006000500040003000200010000FFFFFFFD",
		INIT_5C=>X"FFFEFFFF00010002000300040005000600070008000800090009000A000A000A",
		INIT_5D=>X"FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFD",
		INIT_5E=>X"000500040003000200010000FFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF6",
		INIT_5F=>X"000800080009000A000A000A000B000B000B000A000A000A0009000800070006",
		INIT_60=>X"FFF6FFF6FFF7FFF8FFF9FFFBFFFCFFFDFFFE0000000100020003000400060007",
		INIT_61=>X"FFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF4FFF5FFF5",
		INIT_62=>X"000C000B000B000A000A00090008000700060005000300020001FFFFFFFEFFFD",
		INIT_63=>X"FFFE000000010002000400050006000700080009000A000B000B000C000C000C",
		INIT_64=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFD",
		INIT_65=>X"00060005000400020001FFFFFFFEFFFCFFFBFFFAFFF8FFF7FFF6FFF5FFF4FFF4",
		INIT_66=>X"000A000B000B000C000D000D000D000D000D000D000C000C000B000A00090008",
		INIT_67=>X"FFF4FFF5FFF6FFF7FFF8FFFAFFFBFFFDFFFE0000000100030004000600070008",
		INIT_68=>X"FFFAFFF9FFF7FFF6FFF5FFF4FFF3FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF2FFF3",
		INIT_69=>X"000F000F000E000D000C000B000A000900070006000400020001FFFFFFFDFFFC",
		INIT_6A=>X"FFFE000000020004000500070008000A000B000C000D000E000F000F000F000F",
		INIT_6B=>X"FFEFFFEFFFEFFFEFFFEFFFEFFFF0FFF1FFF2FFF3FFF4FFF6FFF7FFF9FFFBFFFC",
		INIT_6C=>X"00080006000500030001FFFFFFFDFFFBFFF9FFF7FFF6FFF4FFF3FFF2FFF1FFF0",
		INIT_6D=>X"000D000F001000110011001200120012001200110010000F000E000D000C000A",
		INIT_6E=>X"FFEFFFF1FFF2FFF4FFF6FFF8FFFAFFFCFFFE00000003000500070009000A000C",
		INIT_6F=>X"FFF8FFF5FFF3FFF2FFF0FFEFFFEEFFEDFFECFFECFFEBFFEBFFECFFECFFEDFFEE",
		INIT_70=>X"001500150014001300110010000E000C000A0008000500030001FFFEFFFCFFFA",
		INIT_71=>X"FFFE0001000400060009000B000D000F00110012001300140015001600160016",
		INIT_72=>X"FFE7FFE6FFE6FFE6FFE7FFE8FFE9FFEAFFECFFEDFFEFFFF2FFF4FFF6FFF9FFFC",
		INIT_73=>X"000C000A000700040001FFFEFFFBFFF8FFF5FFF2FFF0FFEEFFECFFEAFFE9FFE8",
		INIT_74=>X"00160018001A001B001C001C001D001C001C001B001A0018001600140012000F",
		INIT_75=>X"FFE5FFE8FFEAFFEDFFF1FFF4FFF7FFFBFFFE000200050009000C000F00110014",
		INIT_76=>X"FFF1FFEDFFEAFFE7FFE4FFE2FFE0FFDFFFDEFFDDFFDDFFDEFFDEFFDFFFE1FFE3",
		INIT_77=>X"0028002600240022001F001C001900150011000D000900050001FFFCFFF8FFF4",
		INIT_78=>X"FFFE00040009000D00120016001A001E00210024002600270028002900290029",
		INIT_79=>X"FFCBFFCAFFCAFFCBFFCCFFCEFFD1FFD4FFD7FFDBFFE0FFE4FFE9FFEFFFF4FFF9",
		INIT_7A=>X"001D0016000F00080001FFFAFFF3FFEDFFE7FFE1FFDCFFD8FFD4FFD0FFCEFFCC",
		INIT_7B=>X"003F004300460049004A004B004A0049004700430040003B00360030002A0024",
		INIT_7C=>X"FFAAFFB3FFBEFFC8FFD3FFDEFFE9FFF4FFFE00090012001C0024002C00330039",
		INIT_7D=>X"FFBAFFACFFA1FF97FF8FFF89FF84FF82FF81FF81FF83FF87FF8CFF92FF99FFA1",
		INIT_7E=>X"013E0121010500E900CC00B000940079005F0045002D00160001FFECFFDAFFC9",
		INIT_7F=>X"024802460243023D02340229021D020E01FC01EA01D501BF01A7018E01740159",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_05,
		DOPADOP=>dopadop_05,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_06: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"F00000000000000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF0000000",
		INITP_01=>X"FFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFF",
		INITP_02=>X"000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000000FFFFF",
		INITP_03=>X"00000000000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000",
		INITP_04=>X"FFFFC00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC000",
		INITP_05=>X"FFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFF",
		INITP_06=>X"0000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC00000000000003F",
		INITP_07=>X"000000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC0000000",
		INITP_08=>X"FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFF",
		INITP_09=>X"0000FFFFFFFFFF0000000000FFFFFFFFFF0000000003FFFFFFFFFC0000000003",
		INITP_0A=>X"000000003FFFFFFFFFC000000000FFFFFFFFFF0000000000FFFFFFFFFF000000",
		INITP_0B=>X"FFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0",
		INITP_0C=>X"FFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFF",
		INITP_0D=>X"03FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFF0000000000FFF",
		INITP_0E=>X"000000FFFFFFFFFF0000000003FFFFFFFFFC0000000003FFFFFFFFFC00000000",
		INITP_0F=>X"0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000",
		INIT_00=>X"FFFEFFFF00000000000100020003000400040005000600060007000700070007",
		INIT_01=>X"FFF8FFF8FFF8FFF8FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFD",
		INIT_02=>X"000400040003000200010000FFFFFFFFFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF9",
		INIT_03=>X"0005000500060006000700070007000700080007000700070007000600060005",
		INIT_04=>X"FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFEFFFF000000010001000200030004",
		INIT_05=>X"FFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF9FFF8FFF8FFF8FFF7FFF7FFF8FFF8FFF8",
		INIT_06=>X"00080008000700070007000600060005000400040003000200010000FFFFFFFE",
		INIT_07=>X"FFFEFFFF00000001000200020003000400050005000600060007000700070008",
		INIT_08=>X"FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFD",
		INIT_09=>X"000400040003000200010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFFAFFF9FFF8",
		INIT_0A=>X"0005000600060007000700070008000800080008000700070007000600060005",
		INIT_0B=>X"FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFEFFFF000000010002000300030004",
		INIT_0C=>X"FFFDFFFCFFFCFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF8",
		INIT_0D=>X"00080008000800070007000600060005000400040003000200010000FFFFFFFE",
		INIT_0E=>X"FFFEFFFF00000001000200030004000400050006000600070007000800080008",
		INIT_0F=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFFAFFFBFFFBFFFCFFFD",
		INIT_10=>X"000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8",
		INIT_11=>X"0005000600070007000800080008000800080008000800080007000700060005",
		INIT_12=>X"FFF8FFF8FFF9FFFAFFFAFFFBFFFCFFFDFFFEFFFF000000010002000300040005",
		INIT_13=>X"FFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_14=>X"00090009000800080007000700060005000500040003000200010000FFFFFFFE",
		INIT_15=>X"FFFEFFFF00000001000200030004000500060007000700080008000800090009",
		INIT_16=>X"FFF7FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF9FFF9FFFAFFFBFFFCFFFD",
		INIT_17=>X"000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF7",
		INIT_18=>X"0006000700080008000900090009000900090009000900080008000700070006",
		INIT_19=>X"FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF000000010003000400050005",
		INIT_1A=>X"FFFCFFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF6FFF6FFF6FFF5FFF6FFF6FFF6FFF6",
		INIT_1B=>X"000A000A000900090008000800070006000500040003000200010000FFFFFFFD",
		INIT_1C=>X"FFFEFFFF00010002000300040005000600070008000800090009000A000A000A",
		INIT_1D=>X"FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFD",
		INIT_1E=>X"000500040003000200010000FFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF6",
		INIT_1F=>X"000800080009000A000A000A000B000B000B000A000A000A0009000800070006",
		INIT_20=>X"FFF6FFF6FFF7FFF8FFF9FFFBFFFCFFFDFFFE0000000100020003000400060007",
		INIT_21=>X"FFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF4FFF5FFF5",
		INIT_22=>X"000C000B000B000A000A00090008000700060005000300020001FFFFFFFEFFFD",
		INIT_23=>X"FFFE000000010002000400050006000700080009000A000B000B000C000C000C",
		INIT_24=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFD",
		INIT_25=>X"00060005000400020001FFFFFFFEFFFCFFFBFFFAFFF8FFF7FFF6FFF5FFF4FFF4",
		INIT_26=>X"000A000B000B000C000D000D000D000D000D000D000C000C000B000A00090008",
		INIT_27=>X"FFF4FFF5FFF6FFF7FFF8FFFAFFFBFFFDFFFE0000000100030004000600070008",
		INIT_28=>X"FFFAFFF9FFF7FFF6FFF5FFF4FFF3FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF2FFF3",
		INIT_29=>X"000F000F000E000D000C000B000A000900070006000400020001FFFFFFFDFFFC",
		INIT_2A=>X"FFFE000000020004000500070008000A000B000C000D000E000F000F000F000F",
		INIT_2B=>X"FFEFFFEFFFEFFFEFFFEFFFEFFFF0FFF1FFF2FFF3FFF4FFF6FFF7FFF9FFFBFFFC",
		INIT_2C=>X"00080006000500030001FFFFFFFDFFFBFFF9FFF7FFF6FFF4FFF3FFF2FFF1FFF0",
		INIT_2D=>X"000D000F001000110011001200120012001200110010000F000E000D000C000A",
		INIT_2E=>X"FFEFFFF1FFF2FFF4FFF6FFF8FFFAFFFCFFFE00000003000500070009000A000C",
		INIT_2F=>X"FFF8FFF5FFF3FFF2FFF0FFEFFFEEFFEDFFECFFECFFEBFFEBFFECFFECFFEDFFEE",
		INIT_30=>X"001500150014001300110010000E000C000A0008000500030001FFFEFFFCFFFA",
		INIT_31=>X"FFFE0001000400060009000B000D000F00110012001300140015001600160016",
		INIT_32=>X"FFE7FFE6FFE6FFE6FFE7FFE8FFE9FFEAFFECFFEDFFEFFFF2FFF4FFF6FFF9FFFC",
		INIT_33=>X"000C000A000700040001FFFEFFFBFFF8FFF5FFF2FFF0FFEEFFECFFEAFFE9FFE8",
		INIT_34=>X"00160018001A001B001C001C001D001C001C001B001A0018001600140012000F",
		INIT_35=>X"FFE5FFE8FFEAFFEDFFF1FFF4FFF7FFFBFFFE000200050009000C000F00110014",
		INIT_36=>X"FFF1FFEDFFEAFFE7FFE4FFE2FFE0FFDFFFDEFFDDFFDDFFDEFFDEFFDFFFE1FFE3",
		INIT_37=>X"0028002600240022001F001C001900150011000D000900050001FFFCFFF8FFF4",
		INIT_38=>X"FFFE00040009000D00120016001A001E00210024002600270028002900290029",
		INIT_39=>X"FFCBFFCAFFCAFFCBFFCCFFCEFFD1FFD4FFD7FFDBFFE0FFE4FFE9FFEFFFF4FFF9",
		INIT_3A=>X"001D0016000F00080001FFFAFFF3FFEDFFE7FFE1FFDCFFD8FFD4FFD0FFCEFFCC",
		INIT_3B=>X"003F004300460049004A004B004A0049004700430040003B00360030002A0024",
		INIT_3C=>X"FFAAFFB3FFBEFFC8FFD3FFDEFFE9FFF4FFFE00090012001C0024002C00330039",
		INIT_3D=>X"FFBAFFACFFA1FF97FF8FFF89FF84FF82FF81FF81FF83FF87FF8CFF92FF99FFA1",
		INIT_3E=>X"013E0121010500E900CC00B000940079005F0045002D00160001FFECFFDAFFC9",
		INIT_3F=>X"024802460243023D02340229021D020E01FC01EA01D501BF01A7018E01740159",
		INIT_40=>X"0006000500040003000200010000FFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF8",
		INIT_41=>X"FFFDFFFEFFFF0001000200030004000500060007000700070008000700070007",
		INIT_42=>X"FFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF8FFF8FFF8FFF9FFFAFFFBFFFC",
		INIT_43=>X"000600060007000700080007000700070006000500050003000200010000FFFF",
		INIT_44=>X"FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFBFFFDFFFEFFFF00000002000300040005",
		INIT_45=>X"0006000600050004000300010000FFFFFFFEFFFCFFFBFFFAFFF9FFF9FFF8FFF8",
		INIT_46=>X"FFFCFFFDFFFF0000000100020004000500060006000700070008000800070007",
		INIT_47=>X"FFFEFFFDFFFCFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF8FFF8FFF8FFF9FFFAFFFB",
		INIT_48=>X"000500060007000700080008000800070007000600050004000300020000FFFF",
		INIT_49=>X"FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFDFFFE00000001000200030004",
		INIT_4A=>X"0007000600050004000300020001FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8",
		INIT_4B=>X"FFFCFFFDFFFEFFFF000100020003000400050006000700070008000800080007",
		INIT_4C=>X"FFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF9FFF9FFFA",
		INIT_4D=>X"0005000600070007000800080008000800070007000600050004000200010000",
		INIT_4E=>X"FFF7FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFEFFFF0000000200030004",
		INIT_4F=>X"00080007000600050004000300010000FFFFFFFDFFFCFFFBFFFAFFF9FFF8FFF8",
		INIT_50=>X"FFFBFFFCFFFDFFFF000000010003000400050006000700080008000800080008",
		INIT_51=>X"FFFFFFFEFFFCFFFBFFFAFFF9FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF9FFFA",
		INIT_52=>X"0005000600070008000800080008000800080007000600050004000300020000",
		INIT_53=>X"FFF7FFF7FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFCFFFDFFFE0000000100030004",
		INIT_54=>X"00080008000700060005000400020001FFFFFFFEFFFDFFFBFFFAFFF9FFF8FFF7",
		INIT_55=>X"FFFAFFFBFFFDFFFEFFFF00010002000400050006000700080008000900090009",
		INIT_56=>X"0000FFFEFFFDFFFBFFFAFFF9FFF8FFF7FFF7FFF6FFF6FFF6FFF7FFF7FFF8FFF9",
		INIT_57=>X"0005000600070008000900090009000900090008000700060005000400030001",
		INIT_58=>X"FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF8FFF9FFFBFFFCFFFEFFFF000100020004",
		INIT_59=>X"000900090008000700060005000300020000FFFFFFFDFFFCFFFAFFF9FFF8FFF7",
		INIT_5A=>X"FFF9FFFAFFFCFFFDFFFF00000002000300050006000700080009000900090009",
		INIT_5B=>X"0001FFFFFFFDFFFCFFFAFFF9FFF8FFF7FFF6FFF6FFF5FFF5FFF6FFF6FFF7FFF8",
		INIT_5C=>X"00050006000700080009000A000A000A000A0009000900080006000500040002",
		INIT_5D=>X"FFF6FFF5FFF5FFF5FFF5FFF5FFF6FFF7FFF8FFFAFFFBFFFDFFFE000000020003",
		INIT_5E=>X"000A000A0009000800070006000400030001FFFFFFFEFFFCFFFAFFF9FFF8FFF7",
		INIT_5F=>X"FFF8FFF9FFFAFFFCFFFE00000001000300050006000700090009000A000A000B",
		INIT_60=>X"00010000FFFEFFFCFFFAFFF9FFF7FFF6FFF5FFF5FFF4FFF4FFF4FFF5FFF5FFF6",
		INIT_61=>X"0005000600080009000A000B000B000B000B000B000A00090008000700050003",
		INIT_62=>X"FFF5FFF4FFF4FFF3FFF3FFF4FFF4FFF5FFF7FFF8FFFAFFFBFFFDFFFF00010003",
		INIT_63=>X"000C000C000B000A000900070006000400020000FFFEFFFCFFFAFFF9FFF7FFF6",
		INIT_64=>X"FFF6FFF7FFF9FFFBFFFDFFFF000100030005000600080009000A000B000C000C",
		INIT_65=>X"00030001FFFFFFFCFFFAFFF9FFF7FFF5FFF4FFF3FFF3FFF2FFF2FFF3FFF3FFF4",
		INIT_66=>X"000500060008000A000B000C000D000D000D000D000C000B000A000800070005",
		INIT_67=>X"FFF4FFF2FFF2FFF1FFF1FFF2FFF2FFF3FFF4FFF6FFF8FFFAFFFCFFFE00000002",
		INIT_68=>X"000E000E000E000D000B000A0008000600040001FFFFFFFDFFFBFFF8FFF7FFF5",
		INIT_69=>X"FFF3FFF5FFF7FFF9FFFBFFFD00000002000400070009000A000C000D000E000E",
		INIT_6A=>X"000500020000FFFDFFFBFFF8FFF6FFF4FFF3FFF1FFF0FFF0FFF0FFF0FFF1FFF2",
		INIT_6B=>X"000400070009000B000D000E000F001000100010000F000E000D000B00090007",
		INIT_6C=>X"FFF1FFF0FFEFFFEEFFEEFFEEFFEFFFF0FFF1FFF3FFF5FFF7FFFAFFFCFFFF0002",
		INIT_6D=>X"0012001200110010000F000D000B0008000600030000FFFDFFFBFFF8FFF6FFF3",
		INIT_6E=>X"FFEFFFF1FFF3FFF6FFF8FFFBFFFE000100040007000A000C000E001000110012",
		INIT_6F=>X"000800040001FFFEFFFBFFF8FFF5FFF2FFF0FFEEFFEDFFECFFECFFECFFECFFED",
		INIT_70=>X"00040008000B000E0010001200130014001500150014001300120010000D000A",
		INIT_71=>X"FFEEFFECFFEAFFE9FFE8FFE8FFE9FFEAFFECFFEEFFF0FFF3FFF6FFFAFFFD0001",
		INIT_72=>X"0019001900180017001500130010000D000A00060002FFFEFFFBFFF7FFF4FFF1",
		INIT_73=>X"FFE7FFEAFFEDFFF0FFF4FFF8FFFC000000040008000C000F0012001500170018",
		INIT_74=>X"000D00090004FFFFFFFBFFF6FFF2FFEEFFEBFFE8FFE6FFE4FFE4FFE4FFE4FFE5",
		INIT_75=>X"00040009000E001200160019001C001D001E001F001E001D001B001800150011",
		INIT_76=>X"FFE6FFE3FFE0FFDEFFDDFFDCFFDDFFDEFFE0FFE3FFE7FFEBFFF0FFF5FFFAFFFF",
		INIT_77=>X"002800280028002600240020001C00170012000C00070001FFFBFFF5FFF0FFEB",
		INIT_78=>X"FFD5FFD9FFDDFFE3FFE9FFF0FFF6FFFD0004000B00110017001C002000240026",
		INIT_79=>X"001C0014000B0003FFFBFFF3FFEBFFE4FFDEFFD9FFD5FFD2FFD0FFD0FFD0FFD2",
		INIT_7A=>X"0004000E001800200028002E003300370039003A003900370034002F002A0023",
		INIT_7B=>X"FFCCFFC3FFBDFFB8FFB5FFB4FFB5FFB8FFBCFFC2FFC9FFD2FFDBFFE5FFEFFFFA",
		INIT_7C=>X"0068006900680064005D0055004B003F0032002500170009FFFBFFEDFFE1FFD6",
		INIT_7D=>X"FF66FF75FF86FF9AFFAEFFC4FFDAFFEF00040018002A003B00490055005E0065",
		INIT_7E=>X"00BB008600540026FFFBFFD4FFB2FF94FF7CFF69FF5AFF51FF4DFF4DFF52FF5A",
		INIT_7F=>X"03380334032A0319030202E402C2029A026D023D020901D3019B0163012A00F2",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_06,
		DOPADOP=>dopadop_06,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_07: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFF",
		INITP_01=>X"0000FFFFFFFFFF0000000000FFFFFFFFFF0000000003FFFFFFFFFC0000000003",
		INITP_02=>X"000000003FFFFFFFFFC000000000FFFFFFFFFF0000000000FFFFFFFFFF000000",
		INITP_03=>X"FFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0",
		INITP_04=>X"FFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFF",
		INITP_05=>X"03FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFF0000000000FFF",
		INITP_06=>X"000000FFFFFFFFFF0000000003FFFFFFFFFC0000000003FFFFFFFFFC00000000",
		INITP_07=>X"0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000",
		INITP_08=>X"FFFF00000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC000",
		INITP_09=>X"00003FFFFFFC0000000FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFF",
		INITP_0A=>X"FFFFF0000000FFFFFFF00000003FFFFFFC0000003FFFFFFC0000003FFFFFFC00",
		INITP_0B=>X"000003FFFFFFC0000003FFFFFFC0000000FFFFFFF0000000FFFFFFF0000000FF",
		INITP_0C=>X"FFFFFF0000000FFFFFFF0000000FFFFFFF00000003FFFFFFC0000003FFFFFFC0",
		INITP_0D=>X"0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000000FFFFFFF0000000F",
		INITP_0E=>X"FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFFFFFF00000003FFFFFFC",
		INITP_0F=>X"00000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000000",
		INIT_00=>X"0006000500040003000200010000FFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF8",
		INIT_01=>X"FFFDFFFEFFFF0001000200030004000500060007000700070008000700070007",
		INIT_02=>X"FFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF8FFF8FFF8FFF9FFFAFFFBFFFC",
		INIT_03=>X"000600060007000700080007000700070006000500050003000200010000FFFF",
		INIT_04=>X"FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFBFFFDFFFEFFFF00000002000300040005",
		INIT_05=>X"0006000600050004000300010000FFFFFFFEFFFCFFFBFFFAFFF9FFF9FFF8FFF8",
		INIT_06=>X"FFFCFFFDFFFF0000000100020004000500060006000700070008000800070007",
		INIT_07=>X"FFFEFFFDFFFCFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF8FFF8FFF8FFF9FFFAFFFB",
		INIT_08=>X"000500060007000700080008000800070007000600050004000300020000FFFF",
		INIT_09=>X"FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFDFFFE00000001000200030004",
		INIT_0A=>X"0007000600050004000300020001FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8",
		INIT_0B=>X"FFFCFFFDFFFEFFFF000100020003000400050006000700070008000800080007",
		INIT_0C=>X"FFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF9FFF9FFFA",
		INIT_0D=>X"0005000600070007000800080008000800070007000600050004000200010000",
		INIT_0E=>X"FFF7FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFEFFFF0000000200030004",
		INIT_0F=>X"00080007000600050004000300010000FFFFFFFDFFFCFFFBFFFAFFF9FFF8FFF8",
		INIT_10=>X"FFFBFFFCFFFDFFFF000000010003000400050006000700080008000800080008",
		INIT_11=>X"FFFFFFFEFFFCFFFBFFFAFFF9FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF9FFFA",
		INIT_12=>X"0005000600070008000800080008000800080007000600050004000300020000",
		INIT_13=>X"FFF7FFF7FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFCFFFDFFFE0000000100030004",
		INIT_14=>X"00080008000700060005000400020001FFFFFFFEFFFDFFFBFFFAFFF9FFF8FFF7",
		INIT_15=>X"FFFAFFFBFFFDFFFEFFFF00010002000400050006000700080008000900090009",
		INIT_16=>X"0000FFFEFFFDFFFBFFFAFFF9FFF8FFF7FFF7FFF6FFF6FFF6FFF7FFF7FFF8FFF9",
		INIT_17=>X"0005000600070008000900090009000900090008000700060005000400030001",
		INIT_18=>X"FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF8FFF9FFFBFFFCFFFEFFFF000100020004",
		INIT_19=>X"000900090008000700060005000300020000FFFFFFFDFFFCFFFAFFF9FFF8FFF7",
		INIT_1A=>X"FFF9FFFAFFFCFFFDFFFF00000002000300050006000700080009000900090009",
		INIT_1B=>X"0001FFFFFFFDFFFCFFFAFFF9FFF8FFF7FFF6FFF6FFF5FFF5FFF6FFF6FFF7FFF8",
		INIT_1C=>X"00050006000700080009000A000A000A000A0009000900080006000500040002",
		INIT_1D=>X"FFF6FFF5FFF5FFF5FFF5FFF5FFF6FFF7FFF8FFFAFFFBFFFDFFFE000000020003",
		INIT_1E=>X"000A000A0009000800070006000400030001FFFFFFFEFFFCFFFAFFF9FFF8FFF7",
		INIT_1F=>X"FFF8FFF9FFFAFFFCFFFE00000001000300050006000700090009000A000A000B",
		INIT_20=>X"00010000FFFEFFFCFFFAFFF9FFF7FFF6FFF5FFF5FFF4FFF4FFF4FFF5FFF5FFF6",
		INIT_21=>X"0005000600080009000A000B000B000B000B000B000A00090008000700050003",
		INIT_22=>X"FFF5FFF4FFF4FFF3FFF3FFF4FFF4FFF5FFF7FFF8FFFAFFFBFFFDFFFF00010003",
		INIT_23=>X"000C000C000B000A000900070006000400020000FFFEFFFCFFFAFFF9FFF7FFF6",
		INIT_24=>X"FFF6FFF7FFF9FFFBFFFDFFFF000100030005000600080009000A000B000C000C",
		INIT_25=>X"00030001FFFFFFFCFFFAFFF9FFF7FFF5FFF4FFF3FFF3FFF2FFF2FFF3FFF3FFF4",
		INIT_26=>X"000500060008000A000B000C000D000D000D000D000C000B000A000800070005",
		INIT_27=>X"FFF4FFF2FFF2FFF1FFF1FFF2FFF2FFF3FFF4FFF6FFF8FFFAFFFCFFFE00000002",
		INIT_28=>X"000E000E000E000D000B000A0008000600040001FFFFFFFDFFFBFFF8FFF7FFF5",
		INIT_29=>X"FFF3FFF5FFF7FFF9FFFBFFFD00000002000400070009000A000C000D000E000E",
		INIT_2A=>X"000500020000FFFDFFFBFFF8FFF6FFF4FFF3FFF1FFF0FFF0FFF0FFF0FFF1FFF2",
		INIT_2B=>X"000400070009000B000D000E000F001000100010000F000E000D000B00090007",
		INIT_2C=>X"FFF1FFF0FFEFFFEEFFEEFFEEFFEFFFF0FFF1FFF3FFF5FFF7FFFAFFFCFFFF0002",
		INIT_2D=>X"0012001200110010000F000D000B0008000600030000FFFDFFFBFFF8FFF6FFF3",
		INIT_2E=>X"FFEFFFF1FFF3FFF6FFF8FFFBFFFE000100040007000A000C000E001000110012",
		INIT_2F=>X"000800040001FFFEFFFBFFF8FFF5FFF2FFF0FFEEFFEDFFECFFECFFECFFECFFED",
		INIT_30=>X"00040008000B000E0010001200130014001500150014001300120010000D000A",
		INIT_31=>X"FFEEFFECFFEAFFE9FFE8FFE8FFE9FFEAFFECFFEEFFF0FFF3FFF6FFFAFFFD0001",
		INIT_32=>X"0019001900180017001500130010000D000A00060002FFFEFFFBFFF7FFF4FFF1",
		INIT_33=>X"FFE7FFEAFFEDFFF0FFF4FFF8FFFC000000040008000C000F0012001500170018",
		INIT_34=>X"000D00090004FFFFFFFBFFF6FFF2FFEEFFEBFFE8FFE6FFE4FFE4FFE4FFE4FFE5",
		INIT_35=>X"00040009000E001200160019001C001D001E001F001E001D001B001800150011",
		INIT_36=>X"FFE6FFE3FFE0FFDEFFDDFFDCFFDDFFDEFFE0FFE3FFE7FFEBFFF0FFF5FFFAFFFF",
		INIT_37=>X"002800280028002600240020001C00170012000C00070001FFFBFFF5FFF0FFEB",
		INIT_38=>X"FFD5FFD9FFDDFFE3FFE9FFF0FFF6FFFD0004000B00110017001C002000240026",
		INIT_39=>X"001C0014000B0003FFFBFFF3FFEBFFE4FFDEFFD9FFD5FFD2FFD0FFD0FFD0FFD2",
		INIT_3A=>X"0004000E001800200028002E003300370039003A003900370034002F002A0023",
		INIT_3B=>X"FFCCFFC3FFBDFFB8FFB5FFB4FFB5FFB8FFBCFFC2FFC9FFD2FFDBFFE5FFEFFFFA",
		INIT_3C=>X"0068006900680064005D0055004B003F0032002500170009FFFBFFEDFFE1FFD6",
		INIT_3D=>X"FF66FF75FF86FF9AFFAEFFC4FFDAFFEF00040018002A003B00490055005E0065",
		INIT_3E=>X"00BB008600540026FFFBFFD4FFB2FF94FF7CFF69FF5AFF51FF4DFF4DFF52FF5A",
		INIT_3F=>X"03380334032A0319030202E402C2029A026D023D020901D3019B0163012A00F2",
		INIT_40=>X"FFF8FFF8FFF8FFF8FFF8FFF9FFFBFFFCFFFE0000000100030005000600070007",
		INIT_41=>X"00050006000700070007000700070006000400030001FFFFFFFDFFFCFFFAFFF9",
		INIT_42=>X"FFFDFFFBFFFAFFF9FFF8FFF8FFF8FFF8FFF9FFFAFFFBFFFDFFFE000000020003",
		INIT_43=>X"FFFF00000002000400050006000700070007000700060005000400020001FFFF",
		INIT_44=>X"000300020000FFFEFFFDFFFBFFFAFFF9FFF8FFF7FFF8FFF8FFF9FFFAFFFBFFFD",
		INIT_45=>X"FFF9FFFAFFFCFFFDFFFF00010003000400060007000700080007000700060005",
		INIT_46=>X"0007000700060005000300010000FFFEFFFCFFFBFFF9FFF8FFF8FFF7FFF8FFF8",
		INIT_47=>X"FFF8FFF7FFF8FFF8FFF9FFFBFFFCFFFE00000001000300050006000700070008",
		INIT_48=>X"0006000700080008000700070006000400030001FFFFFFFDFFFCFFFAFFF9FFF8",
		INIT_49=>X"FFFBFFFAFFF9FFF8FFF7FFF7FFF8FFF8FFF9FFFBFFFCFFFE0000000200040005",
		INIT_4A=>X"00010002000400050007000700080008000700070005000400020001FFFFFFFD",
		INIT_4B=>X"00020000FFFEFFFCFFFBFFF9FFF8FFF8FFF7FFF7FFF8FFF9FFFAFFFBFFFDFFFF",
		INIT_4C=>X"FFFAFFFCFFFDFFFF000100030004000600070008000800080007000600050004",
		INIT_4D=>X"000700060005000300020000FFFEFFFCFFFAFFF9FFF8FFF7FFF7FFF7FFF8FFF9",
		INIT_4E=>X"FFF7FFF7FFF8FFF9FFFAFFFCFFFE000000010003000500060007000800080008",
		INIT_4F=>X"000800080008000800070006000500030001FFFFFFFDFFFCFFFAFFF9FFF8FFF7",
		INIT_50=>X"FFF9FFF8FFF7FFF7FFF7FFF7FFF8FFF9FFFBFFFCFFFE00000002000400050007",
		INIT_51=>X"0002000400060007000800080008000800070006000400030001FFFFFFFDFFFB",
		INIT_52=>X"0000FFFEFFFCFFFBFFF9FFF8FFF7FFF7FFF7FFF7FFF8FFF9FFFBFFFDFFFF0001",
		INIT_53=>X"FFFBFFFDFFFF0001000300050006000700080008000800080007000600040002",
		INIT_54=>X"00070005000400020000FFFEFFFCFFFAFFF9FFF7FFF7FFF6FFF7FFF7FFF8FFFA",
		INIT_55=>X"FFF6FFF7FFF8FFFAFFFCFFFE0000000200040005000700080008000900080008",
		INIT_56=>X"00090009000900080007000500030001FFFFFFFDFFFBFFF9FFF8FFF7FFF6FFF6",
		INIT_57=>X"FFF8FFF7FFF6FFF6FFF6FFF7FFF8FFFAFFFCFFFE000000020004000600070008",
		INIT_58=>X"000500060008000900090009000900080006000500030001FFFFFFFDFFFBFFF9",
		INIT_59=>X"FFFEFFFCFFFAFFF8FFF7FFF6FFF6FFF6FFF6FFF7FFF9FFFAFFFCFFFE00010003",
		INIT_5A=>X"FFFDFFFF000100030005000700080009000A0009000900080006000400020000",
		INIT_5B=>X"0006000400020000FFFDFFFBFFF9FFF8FFF6FFF6FFF5FFF5FFF6FFF7FFF9FFFB",
		INIT_5C=>X"FFF6FFF7FFF9FFFBFFFD000000020004000600080009000A000A000A00090008",
		INIT_5D=>X"000A000A00090008000600040001FFFFFFFDFFFBFFF9FFF7FFF6FFF5FFF5FFF5",
		INIT_5E=>X"FFF5FFF5FFF5FFF5FFF6FFF7FFF9FFFBFFFE000000030005000700080009000A",
		INIT_5F=>X"00080009000A000B000B000A00090008000600030001FFFEFFFCFFFAFFF8FFF6",
		INIT_60=>X"FFFBFFF9FFF7FFF6FFF5FFF4FFF4FFF5FFF6FFF8FFFAFFFCFFFE000100030006",
		INIT_61=>X"FFFF0002000400060008000A000B000B000B000A00090007000500030000FFFE",
		INIT_62=>X"000500020000FFFDFFFBFFF8FFF6FFF5FFF4FFF3FFF4FFF4FFF6FFF8FFFAFFFC",
		INIT_63=>X"FFF6FFF8FFFAFFFD00000002000500070009000B000C000C000C000B00090007",
		INIT_64=>X"000C000B0009000700050002FFFFFFFCFFFAFFF7FFF5FFF4FFF3FFF3FFF3FFF4",
		INIT_65=>X"FFF2FFF2FFF3FFF4FFF6FFF8FFFBFFFD0000000300060008000A000C000C000D",
		INIT_66=>X"000B000D000D000D000D000B0009000700040001FFFEFFFBFFF9FFF6FFF4FFF3",
		INIT_67=>X"FFF8FFF5FFF3FFF2FFF1FFF1FFF2FFF4FFF6FFF8FFFBFFFE0001000400070009",
		INIT_68=>X"000200050008000B000C000E000E000E000D000C0009000700040001FFFDFFFA",
		INIT_69=>X"00030000FFFCFFF9FFF6FFF4FFF2FFF1FFF0FFF1FFF2FFF3FFF6FFF8FFFBFFFF",
		INIT_6A=>X"FFF6FFF9FFFC0000000300060009000C000E000F000F000F000E000C00090007",
		INIT_6B=>X"000E000C000A00060003FFFFFFFBFFF8FFF5FFF2FFF0FFEFFFEFFFF0FFF1FFF3",
		INIT_6C=>X"FFEEFFEFFFF0FFF2FFF5FFF9FFFD000100040008000B000E000F001000110010",
		INIT_6D=>X"0011001200120011000F000D000A00060002FFFEFFFAFFF6FFF3FFF1FFEFFFEE",
		INIT_6E=>X"FFF1FFEFFFEDFFECFFECFFEDFFEFFFF2FFF5FFF9FFFD00020006000A000D000F",
		INIT_6F=>X"0008000C000F001200130014001400120010000D000A00050001FFFDFFF8FFF5",
		INIT_70=>X"0000FFFBFFF7FFF2FFEFFFECFFEBFFEAFFEAFFECFFEEFFF1FFF5FFFAFFFE0003",
		INIT_71=>X"FFF5FFFA00000005000A000E0012001400160016001600140011000E000A0005",
		INIT_72=>X"0013000F000A0004FFFFFFF9FFF4FFF0FFECFFE9FFE8FFE7FFE8FFEAFFEDFFF1",
		INIT_73=>X"FFE5FFE8FFEBFFF0FFF5FFFB00010007000C0011001500180019001900180016",
		INIT_74=>X"001D001D001C001900150010000A0003FFFDFFF7FFF1FFECFFE8FFE5FFE4FFE4",
		INIT_75=>X"FFE3FFE0FFDFFFDFFFE1FFE5FFE9FFEFFFF5FFFC0003000A001000150019001C",
		INIT_76=>X"0015001A001F0022002300220020001C00170011000A0002FFFBFFF4FFEDFFE8",
		INIT_77=>X"FFF8FFEFFFE7FFE1FFDCFFD9FFD8FFD9FFDCFFE0FFE6FFEDFFF5FFFD0006000E",
		INIT_78=>X"FFF50000000A0013001C00220027002A002B002A00270021001B0013000A0001",
		INIT_79=>X"00200015000AFFFEFFF2FFE8FFDFFFD7FFD2FFCFFFCEFFD0FFD4FFDAFFE2FFEB",
		INIT_7A=>X"FFC7FFD0FFDBFFE8FFF500030010001C0027002F003500380038003600310029",
		INIT_7B=>X"0051004C00430038002A001A000AFFF9FFEAFFDBFFCFFFC6FFBFFFBCFFBDFFC0",
		INIT_7C=>X"FF98FF95FF98FF9FFFABFFBAFFCDFFE0FFF5000A001D002E003D0048004F0052",
		INIT_7D=>X"0078008900920094008F00830071005B00410026000AFFEFFFD5FFC0FFAEFFA0",
		INIT_7E=>X"FF7BFF48FF24FF0DFF04FF07FF16FF2FFF4FFF76FF9FFFCBFFF5001D00420060",
		INIT_7F=>X"0488047E0462043303F403A7034D02E8027D020E019E012F00C50063000AFFBC",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_07,
		DOPADOP=>dopadop_07,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_08: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFF00000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC000",
		INITP_01=>X"00003FFFFFFC0000000FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFF",
		INITP_02=>X"FFFFF0000000FFFFFFF00000003FFFFFFC0000003FFFFFFC0000003FFFFFFC00",
		INITP_03=>X"000003FFFFFFC0000003FFFFFFC0000000FFFFFFF0000000FFFFFFF0000000FF",
		INITP_04=>X"FFFFFF0000000FFFFFFF0000000FFFFFFF00000003FFFFFFC0000003FFFFFFC0",
		INITP_05=>X"0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000000FFFFFFF0000000F",
		INITP_06=>X"FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFFFFFF00000003FFFFFFC",
		INITP_07=>X"00000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000000",
		INITP_08=>X"FF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00",
		INITP_09=>X"0FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFF",
		INITP_0A=>X"00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF0000",
		INITP_0B=>X"FFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF",
		INITP_0C=>X"000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000F",
		INITP_0D=>X"FF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00",
		INITP_0E=>X"0FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFF",
		INITP_0F=>X"00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF0000",
		INIT_00=>X"FFF8FFF8FFF8FFF8FFF8FFF9FFFBFFFCFFFE0000000100030005000600070007",
		INIT_01=>X"00050006000700070007000700070006000400030001FFFFFFFDFFFCFFFAFFF9",
		INIT_02=>X"FFFDFFFBFFFAFFF9FFF8FFF8FFF8FFF8FFF9FFFAFFFBFFFDFFFE000000020003",
		INIT_03=>X"FFFF00000002000400050006000700070007000700060005000400020001FFFF",
		INIT_04=>X"000300020000FFFEFFFDFFFBFFFAFFF9FFF8FFF7FFF8FFF8FFF9FFFAFFFBFFFD",
		INIT_05=>X"FFF9FFFAFFFCFFFDFFFF00010003000400060007000700080007000700060005",
		INIT_06=>X"0007000700060005000300010000FFFEFFFCFFFBFFF9FFF8FFF8FFF7FFF8FFF8",
		INIT_07=>X"FFF8FFF7FFF8FFF8FFF9FFFBFFFCFFFE00000001000300050006000700070008",
		INIT_08=>X"0006000700080008000700070006000400030001FFFFFFFDFFFCFFFAFFF9FFF8",
		INIT_09=>X"FFFBFFFAFFF9FFF8FFF7FFF7FFF8FFF8FFF9FFFBFFFCFFFE0000000200040005",
		INIT_0A=>X"00010002000400050007000700080008000700070005000400020001FFFFFFFD",
		INIT_0B=>X"00020000FFFEFFFCFFFBFFF9FFF8FFF8FFF7FFF7FFF8FFF9FFFAFFFBFFFDFFFF",
		INIT_0C=>X"FFFAFFFCFFFDFFFF000100030004000600070008000800080007000600050004",
		INIT_0D=>X"000700060005000300020000FFFEFFFCFFFAFFF9FFF8FFF7FFF7FFF7FFF8FFF9",
		INIT_0E=>X"FFF7FFF7FFF8FFF9FFFAFFFCFFFE000000010003000500060007000800080008",
		INIT_0F=>X"000800080008000800070006000500030001FFFFFFFDFFFCFFFAFFF9FFF8FFF7",
		INIT_10=>X"FFF9FFF8FFF7FFF7FFF7FFF7FFF8FFF9FFFBFFFCFFFE00000002000400050007",
		INIT_11=>X"0002000400060007000800080008000800070006000400030001FFFFFFFDFFFB",
		INIT_12=>X"0000FFFEFFFCFFFBFFF9FFF8FFF7FFF7FFF7FFF7FFF8FFF9FFFBFFFDFFFF0001",
		INIT_13=>X"FFFBFFFDFFFF0001000300050006000700080008000800080007000600040002",
		INIT_14=>X"00070005000400020000FFFEFFFCFFFAFFF9FFF7FFF7FFF6FFF7FFF7FFF8FFFA",
		INIT_15=>X"FFF6FFF7FFF8FFFAFFFCFFFE0000000200040005000700080008000900080008",
		INIT_16=>X"00090009000900080007000500030001FFFFFFFDFFFBFFF9FFF8FFF7FFF6FFF6",
		INIT_17=>X"FFF8FFF7FFF6FFF6FFF6FFF7FFF8FFFAFFFCFFFE000000020004000600070008",
		INIT_18=>X"000500060008000900090009000900080006000500030001FFFFFFFDFFFBFFF9",
		INIT_19=>X"FFFEFFFCFFFAFFF8FFF7FFF6FFF6FFF6FFF6FFF7FFF9FFFAFFFCFFFE00010003",
		INIT_1A=>X"FFFDFFFF000100030005000700080009000A0009000900080006000400020000",
		INIT_1B=>X"0006000400020000FFFDFFFBFFF9FFF8FFF6FFF6FFF5FFF5FFF6FFF7FFF9FFFB",
		INIT_1C=>X"FFF6FFF7FFF9FFFBFFFD000000020004000600080009000A000A000A00090008",
		INIT_1D=>X"000A000A00090008000600040001FFFFFFFDFFFBFFF9FFF7FFF6FFF5FFF5FFF5",
		INIT_1E=>X"FFF5FFF5FFF5FFF5FFF6FFF7FFF9FFFBFFFE000000030005000700080009000A",
		INIT_1F=>X"00080009000A000B000B000A00090008000600030001FFFEFFFCFFFAFFF8FFF6",
		INIT_20=>X"FFFBFFF9FFF7FFF6FFF5FFF4FFF4FFF5FFF6FFF8FFFAFFFCFFFE000100030006",
		INIT_21=>X"FFFF0002000400060008000A000B000B000B000A00090007000500030000FFFE",
		INIT_22=>X"000500020000FFFDFFFBFFF8FFF6FFF5FFF4FFF3FFF4FFF4FFF6FFF8FFFAFFFC",
		INIT_23=>X"FFF6FFF8FFFAFFFD00000002000500070009000B000C000C000C000B00090007",
		INIT_24=>X"000C000B0009000700050002FFFFFFFCFFFAFFF7FFF5FFF4FFF3FFF3FFF3FFF4",
		INIT_25=>X"FFF2FFF2FFF3FFF4FFF6FFF8FFFBFFFD0000000300060008000A000C000C000D",
		INIT_26=>X"000B000D000D000D000D000B0009000700040001FFFEFFFBFFF9FFF6FFF4FFF3",
		INIT_27=>X"FFF8FFF5FFF3FFF2FFF1FFF1FFF2FFF4FFF6FFF8FFFBFFFE0001000400070009",
		INIT_28=>X"000200050008000B000C000E000E000E000D000C0009000700040001FFFDFFFA",
		INIT_29=>X"00030000FFFCFFF9FFF6FFF4FFF2FFF1FFF0FFF1FFF2FFF3FFF6FFF8FFFBFFFF",
		INIT_2A=>X"FFF6FFF9FFFC0000000300060009000C000E000F000F000F000E000C00090007",
		INIT_2B=>X"000E000C000A00060003FFFFFFFBFFF8FFF5FFF2FFF0FFEFFFEFFFF0FFF1FFF3",
		INIT_2C=>X"FFEEFFEFFFF0FFF2FFF5FFF9FFFD000100040008000B000E000F001000110010",
		INIT_2D=>X"0011001200120011000F000D000A00060002FFFEFFFAFFF6FFF3FFF1FFEFFFEE",
		INIT_2E=>X"FFF1FFEFFFEDFFECFFECFFEDFFEFFFF2FFF5FFF9FFFD00020006000A000D000F",
		INIT_2F=>X"0008000C000F001200130014001400120010000D000A00050001FFFDFFF8FFF5",
		INIT_30=>X"0000FFFBFFF7FFF2FFEFFFECFFEBFFEAFFEAFFECFFEEFFF1FFF5FFFAFFFE0003",
		INIT_31=>X"FFF5FFFA00000005000A000E0012001400160016001600140011000E000A0005",
		INIT_32=>X"0013000F000A0004FFFFFFF9FFF4FFF0FFECFFE9FFE8FFE7FFE8FFEAFFEDFFF1",
		INIT_33=>X"FFE5FFE8FFEBFFF0FFF5FFFB00010007000C0011001500180019001900180016",
		INIT_34=>X"001D001D001C001900150010000A0003FFFDFFF7FFF1FFECFFE8FFE5FFE4FFE4",
		INIT_35=>X"FFE3FFE0FFDFFFDFFFE1FFE5FFE9FFEFFFF5FFFC0003000A001000150019001C",
		INIT_36=>X"0015001A001F0022002300220020001C00170011000A0002FFFBFFF4FFEDFFE8",
		INIT_37=>X"FFF8FFEFFFE7FFE1FFDCFFD9FFD8FFD9FFDCFFE0FFE6FFEDFFF5FFFD0006000E",
		INIT_38=>X"FFF50000000A0013001C00220027002A002B002A00270021001B0013000A0001",
		INIT_39=>X"00200015000AFFFEFFF2FFE8FFDFFFD7FFD2FFCFFFCEFFD0FFD4FFDAFFE2FFEB",
		INIT_3A=>X"FFC7FFD0FFDBFFE8FFF500030010001C0027002F003500380038003600310029",
		INIT_3B=>X"0051004C00430038002A001A000AFFF9FFEAFFDBFFCFFFC6FFBFFFBCFFBDFFC0",
		INIT_3C=>X"FF98FF95FF98FF9FFFABFFBAFFCDFFE0FFF5000A001D002E003D0048004F0052",
		INIT_3D=>X"0078008900920094008F00830071005B00410026000AFFEFFFD5FFC0FFAEFFA0",
		INIT_3E=>X"FF7BFF48FF24FF0DFF04FF07FF16FF2FFF4FFF76FF9FFFCBFFF5001D00420060",
		INIT_3F=>X"0488047E0462043303F403A7034D02E8027D020E019E012F00C50063000AFFBC",
		INIT_40=>X"00020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF0002000400060007",
		INIT_41=>X"FFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF00020004000600070008000700060004",
		INIT_42=>X"FFF9FFFBFFFDFFFF0002000400060007000800070006000400020000FFFDFFFB",
		INIT_43=>X"0002000400060007000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF8",
		INIT_44=>X"000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF",
		INIT_45=>X"00020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF0002000400060007",
		INIT_46=>X"FFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF00020004000600070008000700060004",
		INIT_47=>X"FFF9FFFAFFFDFFFF0002000400060007000800070006000500020000FFFDFFFB",
		INIT_48=>X"0002000400060007000800070006000500020000FFFDFFFBFFF9FFF8FFF7FFF8",
		INIT_49=>X"000800070006000500020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFAFFFDFFFF",
		INIT_4A=>X"00020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFAFFFDFFFF0002000400060007",
		INIT_4B=>X"FFF9FFF8FFF7FFF7FFF8FFFAFFFCFFFF00020004000600070008000800060005",
		INIT_4C=>X"FFF8FFFAFFFCFFFF0002000400060007000800080007000500030000FFFDFFFB",
		INIT_4D=>X"0002000400060007000800080007000500030000FFFDFFFBFFF9FFF8FFF7FFF7",
		INIT_4E=>X"000800080007000500030000FFFDFFFBFFF9FFF8FFF7FFF7FFF8FFFAFFFCFFFF",
		INIT_4F=>X"00030000FFFDFFFBFFF9FFF8FFF7FFF7FFF8FFFAFFFCFFFF0002000400060007",
		INIT_50=>X"FFF9FFF7FFF7FFF7FFF8FFFAFFFCFFFF00020004000600080008000800070005",
		INIT_51=>X"FFF8FFFAFFFCFFFF0001000400060008000800080007000500030000FFFEFFFB",
		INIT_52=>X"0001000400060008000800080007000500030000FFFEFFFBFFF9FFF7FFF7FFF7",
		INIT_53=>X"000900080007000600030000FFFEFFFBFFF9FFF7FFF7FFF7FFF8FFFAFFFCFFFF",
		INIT_54=>X"00030000FFFEFFFBFFF9FFF7FFF6FFF7FFF8FFF9FFFCFFFF0001000400060008",
		INIT_55=>X"FFF9FFF7FFF6FFF6FFF7FFF9FFFCFFFF00010004000600080009000900070006",
		INIT_56=>X"FFF7FFF9FFFCFFFE0001000400060008000900090008000600030001FFFEFFFB",
		INIT_57=>X"0001000400070008000900090008000600030001FFFEFFFBFFF8FFF7FFF6FFF6",
		INIT_58=>X"000900090008000600040001FFFEFFFBFFF8FFF7FFF6FFF6FFF7FFF9FFFBFFFE",
		INIT_59=>X"00040001FFFEFFFBFFF8FFF7FFF6FFF6FFF7FFF9FFFBFFFE0001000400070008",
		INIT_5A=>X"FFF8FFF6FFF5FFF6FFF7FFF9FFFBFFFE00010004000700090009000900080006",
		INIT_5B=>X"FFF6FFF8FFFBFFFE0001000400070009000A000A0008000700040001FFFEFFFB",
		INIT_5C=>X"0001000400070009000A000A0009000700040001FFFEFFFBFFF8FFF6FFF5FFF5",
		INIT_5D=>X"000A000A0009000700040001FFFEFFFBFFF8FFF6FFF5FFF5FFF6FFF8FFFBFFFE",
		INIT_5E=>X"00040001FFFEFFFAFFF8FFF6FFF5FFF5FFF6FFF8FFFBFFFE0001000500070009",
		INIT_5F=>X"FFF8FFF5FFF4FFF4FFF5FFF8FFFAFFFE0001000500070009000A000A00090007",
		INIT_60=>X"FFF5FFF7FFFAFFFE000100050008000A000B000B000A000800050001FFFEFFFA",
		INIT_61=>X"000100050008000A000B000B000A000800050001FFFEFFFAFFF7FFF5FFF4FFF4",
		INIT_62=>X"000C000C000A000800050002FFFEFFFAFFF7FFF5FFF4FFF4FFF5FFF7FFFAFFFE",
		INIT_63=>X"00050002FFFEFFFAFFF7FFF4FFF3FFF3FFF4FFF7FFFAFFFD000100050008000A",
		INIT_64=>X"FFF7FFF4FFF3FFF3FFF4FFF6FFF9FFFD000100050008000B000C000C000B0009",
		INIT_65=>X"FFF3FFF6FFF9FFFD000100050009000B000C000D000B000900060002FFFEFFFA",
		INIT_66=>X"000100050009000C000D000D000C000900060002FFFEFFFAFFF6FFF4FFF2FFF2",
		INIT_67=>X"000E000E000D000A00060002FFFEFFFAFFF6FFF3FFF2FFF2FFF3FFF5FFF9FFFD",
		INIT_68=>X"00070002FFFEFFF9FFF5FFF3FFF1FFF1FFF2FFF5FFF8FFFD000100060009000C",
		INIT_69=>X"FFF5FFF2FFF0FFF0FFF1FFF4FFF8FFFC00010006000A000D000E000E000D000B",
		INIT_6A=>X"FFF1FFF3FFF7FFFC00010006000A000D000F000F000E000B00070003FFFEFFF9",
		INIT_6B=>X"00010006000B000E00100010000F000C00080003FFFEFFF9FFF5FFF1FFF0FFEF",
		INIT_6C=>X"001100110010000D00080003FFFEFFF9FFF4FFF1FFEFFFEEFFF0FFF3FFF7FFFC",
		INIT_6D=>X"00090004FFFEFFF8FFF3FFF0FFEEFFEDFFEFFFF2FFF6FFFC00010007000B000F",
		INIT_6E=>X"FFF3FFEFFFECFFECFFEEFFF1FFF6FFFB00010007000C0010001200120011000E",
		INIT_6F=>X"FFECFFF0FFF5FFFB00010007000D0011001300140012000F000A0004FFFEFFF8",
		INIT_70=>X"00010008000E00120015001500140010000B0005FFFEFFF7FFF2FFEDFFEBFFEB",
		INIT_71=>X"0017001700150011000C0005FFFEFFF7FFF1FFECFFE9FFE9FFEBFFEEFFF4FFFA",
		INIT_72=>X"000D0006FFFEFFF6FFEFFFEAFFE7FFE7FFE9FFEDFFF3FFFA00010008000F0014",
		INIT_73=>X"FFEEFFE8FFE5FFE4FFE6FFEBFFF1FFF900010009001000160019001900170013",
		INIT_74=>X"FFE4FFE8FFEFFFF80001000A00120018001B001C001A0015000F0007FFFEFFF5",
		INIT_75=>X"0001000B0014001B001F001F001D001800110008FFFEFFF4FFECFFE6FFE2FFE1",
		INIT_76=>X"002300240021001B00130009FFFEFFF3FFEAFFE3FFDFFFDEFFE0FFE5FFEDFFF7",
		INIT_77=>X"0016000BFFFEFFF2FFE7FFDFFFDAFFD9FFDBFFE1FFEAFFF50001000D0017001E",
		INIT_78=>X"FFE3FFD9FFD3FFD2FFD5FFDCFFE7FFF30001000E001A00230028002900270020",
		INIT_79=>X"FFCCFFD5FFE1FFF100010011001F002A00300031002E0026001B000DFFFEFFEF",
		INIT_7A=>X"0001001500260033003B003D0039002F00210010FFFEFFECFFDDFFD1FFCAFFC8",
		INIT_7B=>X"004E0050004A003E002B0015FFFEFFE7FFD4FFC5FFBCFFBAFFBFFFCAFFD9FFED",
		INIT_7C=>X"003E001FFFFEFFDEFFC3FFAFFFA3FFA1FFA7FFB6FFCCFFE60001001B00320044",
		INIT_7D=>X"FF9EFF7FFF6DFF6AFF76FF8EFFB0FFD800010028004A006300710073006B0058",
		INIT_7E=>X"FECAFF08FF56FFAC0001004E008C00B800CF00D000BE009B006C0036FFFEFFCA",
		INIT_7F=>X"0668064D05FE057F04D80413033A0259017D00B1FFFEFF6BFEFFFEBAFE9DFEA4",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_08,
		DOPADOP=>dopadop_08,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_09: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00",
		INITP_01=>X"0FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFF",
		INITP_02=>X"00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF0000",
		INITP_03=>X"FFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF",
		INITP_04=>X"000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000F",
		INITP_05=>X"FF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00",
		INITP_06=>X"0FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFF",
		INITP_07=>X"00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF0000",
		INITP_08=>X"FF0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC000FFFF0003FFF0003F",
		INITP_09=>X"FC000FFFC0003FFF0003FFF0003FFF0003FFFC000FFFC000FFFC000FFFC000FF",
		INITP_0A=>X"FC000FFFC000FFFC000FFFF0003FFF0003FFF0003FFF0003FFFC000FFFC000FF",
		INITP_0B=>X"F0003FFFC000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF0003FFF0000FF",
		INITP_0C=>X"F0003FFF0003FFF0000FFFC000FFFC000FFFC000FFFC0003FFF0003FFF0003FF",
		INITP_0D=>X"C0003FFF0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC000FFFF0003FF",
		INITP_0E=>X"C000FFFC000FFFC0003FFF0003FFF0003FFF0003FFFC000FFFC000FFFC000FFF",
		INITP_0F=>X"0000FFFC000FFFC000FFFC000FFFF0003FFF0003FFF0003FFF0000FFFC000FFF",
		INIT_00=>X"00020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF0002000400060007",
		INIT_01=>X"FFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF00020004000600070008000700060004",
		INIT_02=>X"FFF9FFFBFFFDFFFF0002000400060007000800070006000400020000FFFDFFFB",
		INIT_03=>X"0002000400060007000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF8",
		INIT_04=>X"000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF",
		INIT_05=>X"00020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF0002000400060007",
		INIT_06=>X"FFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF00020004000600070008000700060004",
		INIT_07=>X"FFF9FFFAFFFDFFFF0002000400060007000800070006000500020000FFFDFFFB",
		INIT_08=>X"0002000400060007000800070006000500020000FFFDFFFBFFF9FFF8FFF7FFF8",
		INIT_09=>X"000800070006000500020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFAFFFDFFFF",
		INIT_0A=>X"00020000FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFAFFFDFFFF0002000400060007",
		INIT_0B=>X"FFF9FFF8FFF7FFF7FFF8FFFAFFFCFFFF00020004000600070008000800060005",
		INIT_0C=>X"FFF8FFFAFFFCFFFF0002000400060007000800080007000500030000FFFDFFFB",
		INIT_0D=>X"0002000400060007000800080007000500030000FFFDFFFBFFF9FFF8FFF7FFF7",
		INIT_0E=>X"000800080007000500030000FFFDFFFBFFF9FFF8FFF7FFF7FFF8FFFAFFFCFFFF",
		INIT_0F=>X"00030000FFFDFFFBFFF9FFF8FFF7FFF7FFF8FFFAFFFCFFFF0002000400060007",
		INIT_10=>X"FFF9FFF7FFF7FFF7FFF8FFFAFFFCFFFF00020004000600080008000800070005",
		INIT_11=>X"FFF8FFFAFFFCFFFF0001000400060008000800080007000500030000FFFEFFFB",
		INIT_12=>X"0001000400060008000800080007000500030000FFFEFFFBFFF9FFF7FFF7FFF7",
		INIT_13=>X"000900080007000600030000FFFEFFFBFFF9FFF7FFF7FFF7FFF8FFFAFFFCFFFF",
		INIT_14=>X"00030000FFFEFFFBFFF9FFF7FFF6FFF7FFF8FFF9FFFCFFFF0001000400060008",
		INIT_15=>X"FFF9FFF7FFF6FFF6FFF7FFF9FFFCFFFF00010004000600080009000900070006",
		INIT_16=>X"FFF7FFF9FFFCFFFE0001000400060008000900090008000600030001FFFEFFFB",
		INIT_17=>X"0001000400070008000900090008000600030001FFFEFFFBFFF8FFF7FFF6FFF6",
		INIT_18=>X"000900090008000600040001FFFEFFFBFFF8FFF7FFF6FFF6FFF7FFF9FFFBFFFE",
		INIT_19=>X"00040001FFFEFFFBFFF8FFF7FFF6FFF6FFF7FFF9FFFBFFFE0001000400070008",
		INIT_1A=>X"FFF8FFF6FFF5FFF6FFF7FFF9FFFBFFFE00010004000700090009000900080006",
		INIT_1B=>X"FFF6FFF8FFFBFFFE0001000400070009000A000A0008000700040001FFFEFFFB",
		INIT_1C=>X"0001000400070009000A000A0009000700040001FFFEFFFBFFF8FFF6FFF5FFF5",
		INIT_1D=>X"000A000A0009000700040001FFFEFFFBFFF8FFF6FFF5FFF5FFF6FFF8FFFBFFFE",
		INIT_1E=>X"00040001FFFEFFFAFFF8FFF6FFF5FFF5FFF6FFF8FFFBFFFE0001000500070009",
		INIT_1F=>X"FFF8FFF5FFF4FFF4FFF5FFF8FFFAFFFE0001000500070009000A000A00090007",
		INIT_20=>X"FFF5FFF7FFFAFFFE000100050008000A000B000B000A000800050001FFFEFFFA",
		INIT_21=>X"000100050008000A000B000B000A000800050001FFFEFFFAFFF7FFF5FFF4FFF4",
		INIT_22=>X"000C000C000A000800050002FFFEFFFAFFF7FFF5FFF4FFF4FFF5FFF7FFFAFFFE",
		INIT_23=>X"00050002FFFEFFFAFFF7FFF4FFF3FFF3FFF4FFF7FFFAFFFD000100050008000A",
		INIT_24=>X"FFF7FFF4FFF3FFF3FFF4FFF6FFF9FFFD000100050008000B000C000C000B0009",
		INIT_25=>X"FFF3FFF6FFF9FFFD000100050009000B000C000D000B000900060002FFFEFFFA",
		INIT_26=>X"000100050009000C000D000D000C000900060002FFFEFFFAFFF6FFF4FFF2FFF2",
		INIT_27=>X"000E000E000D000A00060002FFFEFFFAFFF6FFF3FFF2FFF2FFF3FFF5FFF9FFFD",
		INIT_28=>X"00070002FFFEFFF9FFF5FFF3FFF1FFF1FFF2FFF5FFF8FFFD000100060009000C",
		INIT_29=>X"FFF5FFF2FFF0FFF0FFF1FFF4FFF8FFFC00010006000A000D000E000E000D000B",
		INIT_2A=>X"FFF1FFF3FFF7FFFC00010006000A000D000F000F000E000B00070003FFFEFFF9",
		INIT_2B=>X"00010006000B000E00100010000F000C00080003FFFEFFF9FFF5FFF1FFF0FFEF",
		INIT_2C=>X"001100110010000D00080003FFFEFFF9FFF4FFF1FFEFFFEEFFF0FFF3FFF7FFFC",
		INIT_2D=>X"00090004FFFEFFF8FFF3FFF0FFEEFFEDFFEFFFF2FFF6FFFC00010007000B000F",
		INIT_2E=>X"FFF3FFEFFFECFFECFFEEFFF1FFF6FFFB00010007000C0010001200120011000E",
		INIT_2F=>X"FFECFFF0FFF5FFFB00010007000D0011001300140012000F000A0004FFFEFFF8",
		INIT_30=>X"00010008000E00120015001500140010000B0005FFFEFFF7FFF2FFEDFFEBFFEB",
		INIT_31=>X"0017001700150011000C0005FFFEFFF7FFF1FFECFFE9FFE9FFEBFFEEFFF4FFFA",
		INIT_32=>X"000D0006FFFEFFF6FFEFFFEAFFE7FFE7FFE9FFEDFFF3FFFA00010008000F0014",
		INIT_33=>X"FFEEFFE8FFE5FFE4FFE6FFEBFFF1FFF900010009001000160019001900170013",
		INIT_34=>X"FFE4FFE8FFEFFFF80001000A00120018001B001C001A0015000F0007FFFEFFF5",
		INIT_35=>X"0001000B0014001B001F001F001D001800110008FFFEFFF4FFECFFE6FFE2FFE1",
		INIT_36=>X"002300240021001B00130009FFFEFFF3FFEAFFE3FFDFFFDEFFE0FFE5FFEDFFF7",
		INIT_37=>X"0016000BFFFEFFF2FFE7FFDFFFDAFFD9FFDBFFE1FFEAFFF50001000D0017001E",
		INIT_38=>X"FFE3FFD9FFD3FFD2FFD5FFDCFFE7FFF30001000E001A00230028002900270020",
		INIT_39=>X"FFCCFFD5FFE1FFF100010011001F002A00300031002E0026001B000DFFFEFFEF",
		INIT_3A=>X"0001001500260033003B003D0039002F00210010FFFEFFECFFDDFFD1FFCAFFC8",
		INIT_3B=>X"004E0050004A003E002B0015FFFEFFE7FFD4FFC5FFBCFFBAFFBFFFCAFFD9FFED",
		INIT_3C=>X"003E001FFFFEFFDEFFC3FFAFFFA3FFA1FFA7FFB6FFCCFFE60001001B00320044",
		INIT_3D=>X"FF9EFF7FFF6DFF6AFF76FF8EFFB0FFD800010028004A006300710073006B0058",
		INIT_3E=>X"FECAFF08FF56FFAC0001004E008C00B800CF00D000BE009B006C0036FFFEFFCA",
		INIT_3F=>X"0668064D05FE057F04D80413033A0259017D00B1FFFEFF6BFEFFFEBAFE9DFEA4",
		INIT_40=>X"FFFAFFF8FFF8FFF9FFFBFFFE0002000500070007000700040001FFFEFFFAFFF8",
		INIT_41=>X"FFFFFFFCFFF9FFF8FFF8FFF9FFFCFFFF0003000600070007000600030000FFFD",
		INIT_42=>X"00050002FFFEFFFBFFF9FFF8FFF8FFFAFFFD0000000400060007000700050003",
		INIT_43=>X"0008000600040001FFFDFFFAFFF8FFF7FFF8FFFBFFFE00010004000700080007",
		INIT_44=>X"000600070007000600030000FFFCFFF9FFF8FFF8FFF9FFFBFFFF000200050007",
		INIT_45=>X"0001000400060008000700050002FFFFFFFBFFF9FFF8FFF8FFF9FFFC00000003",
		INIT_46=>X"FFFBFFFE0002000500070008000700050001FFFEFFFBFFF8FFF7FFF8FFFAFFFD",
		INIT_47=>X"FFF8FFF9FFFCFFFF0003000500070008000600040000FFFDFFFAFFF8FFF7FFF8",
		INIT_48=>X"FFF9FFF7FFF8FFFAFFFD0000000300060008000700060003FFFFFFFCFFF9FFF8",
		INIT_49=>X"FFFDFFFAFFF8FFF7FFF8FFFAFFFD0001000400070008000700050002FFFEFFFB",
		INIT_4A=>X"00040000FFFDFFFAFFF8FFF7FFF8FFFBFFFE0002000500070008000700040001",
		INIT_4B=>X"000800060003FFFFFFFCFFF9FFF7FFF7FFF9FFFCFFFF00030006000800080006",
		INIT_4C=>X"00070008000700050002FFFEFFFBFFF8FFF7FFF8FFFAFFFD0000000400060008",
		INIT_4D=>X"0002000500070008000700040001FFFDFFFAFFF8FFF7FFF8FFFAFFFE00010005",
		INIT_4E=>X"FFFC00000003000600080008000600030000FFFCFFF9FFF7FFF7FFF8FFFBFFFF",
		INIT_4F=>X"FFF8FFFAFFFD0001000400070008000800060003FFFFFFFBFFF8FFF7FFF7FFF9",
		INIT_50=>X"FFF7FFF7FFF8FFFAFFFE0002000500070008000700050002FFFEFFFAFFF8FFF7",
		INIT_51=>X"FFFCFFF9FFF7FFF7FFF8FFFBFFFF0003000600080008000700040001FFFDFFF9",
		INIT_52=>X"0002FFFEFFFBFFF8FFF7FFF7FFF9FFFC0000000400070008000800060003FFFF",
		INIT_53=>X"000800050001FFFDFFFAFFF7FFF6FFF7FFFAFFFD000100050007000800080006",
		INIT_54=>X"00080009000700040000FFFCFFF9FFF7FFF6FFF8FFFBFFFE0002000600080009",
		INIT_55=>X"000400070009000800060003FFFFFFFBFFF8FFF6FFF7FFF8FFFBFFFF00030006",
		INIT_56=>X"FFFD0002000500080009000800060002FFFEFFFAFFF7FFF6FFF7FFF9FFFC0000",
		INIT_57=>X"FFF8FFFBFFFF0003000600080009000800050001FFFDFFF9FFF7FFF6FFF7FFFA",
		INIT_58=>X"FFF6FFF6FFF8FFFC00000004000700090009000700040000FFFCFFF8FFF6FFF6",
		INIT_59=>X"FFFAFFF7FFF6FFF6FFF9FFFD0001000500080009000900070003FFFFFFFBFFF7",
		INIT_5A=>X"0001FFFCFFF9FFF6FFF5FFF7FFFAFFFE000200060009000A000900060002FFFE",
		INIT_5B=>X"000800040000FFFBFFF8FFF6FFF5FFF7FFFBFFFF000300070009000A00080005",
		INIT_5C=>X"000A000900070003FFFEFFFAFFF7FFF5FFF6FFF8FFFC000000040008000A000A",
		INIT_5D=>X"00070009000A000900060002FFFDFFF9FFF6FFF5FFF6FFF9FFFD000100060009",
		INIT_5E=>X"FFFF00040008000A000A000900050000FFFCFFF8FFF5FFF5FFF6FFFAFFFE0003",
		INIT_5F=>X"FFF8FFFC000100050009000B000A00080004FFFFFFFAFFF7FFF5FFF5FFF7FFFB",
		INIT_60=>X"FFF4FFF5FFF8FFFD00020007000A000B000A00070003FFFEFFF9FFF6FFF4FFF5",
		INIT_61=>X"FFF7FFF4FFF4FFF6FFF9FFFE00030008000B000B000A00060001FFFCFFF8FFF5",
		INIT_62=>X"FFFFFFF9FFF6FFF4FFF4FFF6FFFA000000050009000B000B000900050000FFFB",
		INIT_63=>X"00080003FFFDFFF8FFF4FFF3FFF4FFF7FFFC00010006000A000C000B00080004",
		INIT_64=>X"000C000A00060001FFFCFFF7FFF4FFF3FFF4FFF8FFFD00030008000B000C000B",
		INIT_65=>X"000A000D000C000A00050000FFFAFFF5FFF3FFF3FFF5FFF9FFFF00040009000C",
		INIT_66=>X"00020007000C000D000C00090004FFFEFFF8FFF4FFF2FFF3FFF6FFFA00000006",
		INIT_67=>X"FFF8FFFD00040009000D000E000C00080002FFFCFFF7FFF3FFF1FFF3FFF6FFFC",
		INIT_68=>X"FFF1FFF4FFF9FFFF0005000B000E000E000C00070001FFFAFFF5FFF2FFF1FFF3",
		INIT_69=>X"FFF2FFF0FFF1FFF5FFFA00010007000C000F000E000B0006FFFFFFF9FFF4FFF1",
		INIT_6A=>X"FFFBFFF5FFF1FFEFFFF1FFF6FFFC00030009000E000F000E000A0004FFFDFFF7",
		INIT_6B=>X"00080000FFF9FFF3FFEFFFEFFFF2FFF7FFFE0005000B000F0010000E00090002",
		INIT_6C=>X"0010000C0006FFFEFFF7FFF1FFEEFFEFFFF2FFF800000007000D00100010000D",
		INIT_6D=>X"001000120010000B0004FFFCFFF5FFEFFFEDFFEFFFF3FFFA00020009000F0011",
		INIT_6E=>X"0007000E001200130010000A0002FFFAFFF2FFEEFFECFFEFFFF4FFFC0004000B",
		INIT_6F=>X"FFF800000009001000140013000F00080000FFF7FFF0FFECFFECFFEFFFF6FFFE",
		INIT_70=>X"FFEBFFF1FFFA0003000C001200150014000F0007FFFDFFF4FFEEFFEBFFEBFFF0",
		INIT_71=>X"FFE9FFE8FFEBFFF2FFFC0006000F001500160014000D0004FFFAFFF2FFEBFFE9",
		INIT_72=>X"FFF4FFECFFE7FFE7FFECFFF4FFFF00090012001700180014000C0002FFF7FFEF",
		INIT_73=>X"0008FFFCFFF0FFE8FFE5FFE6FFECFFF60002000D0015001900190013000AFFFF",
		INIT_74=>X"001A00110005FFF8FFECFFE5FFE2FFE6FFEEFFF9000500110018001B00190012",
		INIT_75=>X"001F0020001A000F0001FFF4FFE8FFE1FFE0FFE5FFEFFFFC00090015001C001E",
		INIT_76=>X"0013001E002300220019000CFFFDFFEFFFE3FFDEFFDEFFE5FFF10000000E0019",
		INIT_77=>X"FFF80009001900240027002300190009FFF8FFE9FFDEFFDAFFDDFFE6FFF40004",
		INIT_78=>X"FFD9FFE9FFFC00100020002A002C002500170005FFF3FFE3FFD8FFD6FFDBFFE7",
		INIT_79=>X"FFCAFFCCFFD8FFEB00020018002800310030002600150000FFECFFDBFFD2FFD1",
		INIT_7A=>X"FFD7FFC6FFC0FFC6FFD7FFEF000900220033003A003600280012FFFAFFE3FFD2",
		INIT_7B=>X"0008FFE5FFC8FFB6FFB3FFBEFFD5FFF40014002F00400045003D0029000EFFF1",
		INIT_7C=>X"0052002BFFFDFFD2FFB1FFA0FFA1FFB4FFD5FFFC00230042005300540045002A",
		INIT_7D=>X"00A200920067002BFFEBFFB2FF8AFF7AFF84FFA4FFD40009003B005F006F006A",
		INIT_7E=>X"00E0011E012100EF0097002CFFC2FF6DFF3AFF2FFF4BFF86FFD3002300680094",
		INIT_7F=>X"08F808AE07DA06940500034A01A0002CFF0DFE58FE0FFE29FE92FF2AFFD3006D",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_09,
		DOPADOP=>dopadop_09,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_10: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FF0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC000FFFF0003FFF0003F",
		INITP_01=>X"FC000FFFC0003FFF0003FFF0003FFF0003FFFC000FFFC000FFFC000FFFC000FF",
		INITP_02=>X"FC000FFFC000FFFC000FFFF0003FFF0003FFF0003FFF0003FFFC000FFFC000FF",
		INITP_03=>X"F0003FFFC000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF0003FFF0000FF",
		INITP_04=>X"F0003FFF0003FFF0000FFFC000FFFC000FFFC000FFFC0003FFF0003FFF0003FF",
		INITP_05=>X"C0003FFF0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC000FFFF0003FF",
		INITP_06=>X"C000FFFC000FFFC0003FFF0003FFF0003FFF0003FFFC000FFFC000FFFC000FFF",
		INITP_07=>X"0000FFFC000FFFC000FFFC000FFFF0003FFF0003FFF0003FFF0000FFFC000FFF",
		INITP_08=>X"00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF003FFC00FFC00FFC00F",
		INITP_09=>X"FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FF000FFC00FFC00FFC",
		INITP_0A=>X"C00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FF000FFC00FFC00",
		INITP_0B=>X"0FFC00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF003FF000FFC00FF",
		INITP_0C=>X"FC00FFC00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF003FFC00FFC0",
		INITP_0D=>X"00FFC00FFC00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF003FFC00F",
		INITP_0E=>X"FFC00FFC00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FF000FFC",
		INITP_0F=>X"000FFC00FFC00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FF000",
		INIT_00=>X"FFFAFFF8FFF8FFF9FFFBFFFE0002000500070007000700040001FFFEFFFAFFF8",
		INIT_01=>X"FFFFFFFCFFF9FFF8FFF8FFF9FFFCFFFF0003000600070007000600030000FFFD",
		INIT_02=>X"00050002FFFEFFFBFFF9FFF8FFF8FFFAFFFD0000000400060007000700050003",
		INIT_03=>X"0008000600040001FFFDFFFAFFF8FFF7FFF8FFFBFFFE00010004000700080007",
		INIT_04=>X"000600070007000600030000FFFCFFF9FFF8FFF8FFF9FFFBFFFF000200050007",
		INIT_05=>X"0001000400060008000700050002FFFFFFFBFFF9FFF8FFF8FFF9FFFC00000003",
		INIT_06=>X"FFFBFFFE0002000500070008000700050001FFFEFFFBFFF8FFF7FFF8FFFAFFFD",
		INIT_07=>X"FFF8FFF9FFFCFFFF0003000500070008000600040000FFFDFFFAFFF8FFF7FFF8",
		INIT_08=>X"FFF9FFF7FFF8FFFAFFFD0000000300060008000700060003FFFFFFFCFFF9FFF8",
		INIT_09=>X"FFFDFFFAFFF8FFF7FFF8FFFAFFFD0001000400070008000700050002FFFEFFFB",
		INIT_0A=>X"00040000FFFDFFFAFFF8FFF7FFF8FFFBFFFE0002000500070008000700040001",
		INIT_0B=>X"000800060003FFFFFFFCFFF9FFF7FFF7FFF9FFFCFFFF00030006000800080006",
		INIT_0C=>X"00070008000700050002FFFEFFFBFFF8FFF7FFF8FFFAFFFD0000000400060008",
		INIT_0D=>X"0002000500070008000700040001FFFDFFFAFFF8FFF7FFF8FFFAFFFE00010005",
		INIT_0E=>X"FFFC00000003000600080008000600030000FFFCFFF9FFF7FFF7FFF8FFFBFFFF",
		INIT_0F=>X"FFF8FFFAFFFD0001000400070008000800060003FFFFFFFBFFF8FFF7FFF7FFF9",
		INIT_10=>X"FFF7FFF7FFF8FFFAFFFE0002000500070008000700050002FFFEFFFAFFF8FFF7",
		INIT_11=>X"FFFCFFF9FFF7FFF7FFF8FFFBFFFF0003000600080008000700040001FFFDFFF9",
		INIT_12=>X"0002FFFEFFFBFFF8FFF7FFF7FFF9FFFC0000000400070008000800060003FFFF",
		INIT_13=>X"000800050001FFFDFFFAFFF7FFF6FFF7FFFAFFFD000100050007000800080006",
		INIT_14=>X"00080009000700040000FFFCFFF9FFF7FFF6FFF8FFFBFFFE0002000600080009",
		INIT_15=>X"000400070009000800060003FFFFFFFBFFF8FFF6FFF7FFF8FFFBFFFF00030006",
		INIT_16=>X"FFFD0002000500080009000800060002FFFEFFFAFFF7FFF6FFF7FFF9FFFC0000",
		INIT_17=>X"FFF8FFFBFFFF0003000600080009000800050001FFFDFFF9FFF7FFF6FFF7FFFA",
		INIT_18=>X"FFF6FFF6FFF8FFFC00000004000700090009000700040000FFFCFFF8FFF6FFF6",
		INIT_19=>X"FFFAFFF7FFF6FFF6FFF9FFFD0001000500080009000900070003FFFFFFFBFFF7",
		INIT_1A=>X"0001FFFCFFF9FFF6FFF5FFF7FFFAFFFE000200060009000A000900060002FFFE",
		INIT_1B=>X"000800040000FFFBFFF8FFF6FFF5FFF7FFFBFFFF000300070009000A00080005",
		INIT_1C=>X"000A000900070003FFFEFFFAFFF7FFF5FFF6FFF8FFFC000000040008000A000A",
		INIT_1D=>X"00070009000A000900060002FFFDFFF9FFF6FFF5FFF6FFF9FFFD000100060009",
		INIT_1E=>X"FFFF00040008000A000A000900050000FFFCFFF8FFF5FFF5FFF6FFFAFFFE0003",
		INIT_1F=>X"FFF8FFFC000100050009000B000A00080004FFFFFFFAFFF7FFF5FFF5FFF7FFFB",
		INIT_20=>X"FFF4FFF5FFF8FFFD00020007000A000B000A00070003FFFEFFF9FFF6FFF4FFF5",
		INIT_21=>X"FFF7FFF4FFF4FFF6FFF9FFFE00030008000B000B000A00060001FFFCFFF8FFF5",
		INIT_22=>X"FFFFFFF9FFF6FFF4FFF4FFF6FFFA000000050009000B000B000900050000FFFB",
		INIT_23=>X"00080003FFFDFFF8FFF4FFF3FFF4FFF7FFFC00010006000A000C000B00080004",
		INIT_24=>X"000C000A00060001FFFCFFF7FFF4FFF3FFF4FFF8FFFD00030008000B000C000B",
		INIT_25=>X"000A000D000C000A00050000FFFAFFF5FFF3FFF3FFF5FFF9FFFF00040009000C",
		INIT_26=>X"00020007000C000D000C00090004FFFEFFF8FFF4FFF2FFF3FFF6FFFA00000006",
		INIT_27=>X"FFF8FFFD00040009000D000E000C00080002FFFCFFF7FFF3FFF1FFF3FFF6FFFC",
		INIT_28=>X"FFF1FFF4FFF9FFFF0005000B000E000E000C00070001FFFAFFF5FFF2FFF1FFF3",
		INIT_29=>X"FFF2FFF0FFF1FFF5FFFA00010007000C000F000E000B0006FFFFFFF9FFF4FFF1",
		INIT_2A=>X"FFFBFFF5FFF1FFEFFFF1FFF6FFFC00030009000E000F000E000A0004FFFDFFF7",
		INIT_2B=>X"00080000FFF9FFF3FFEFFFEFFFF2FFF7FFFE0005000B000F0010000E00090002",
		INIT_2C=>X"0010000C0006FFFEFFF7FFF1FFEEFFEFFFF2FFF800000007000D00100010000D",
		INIT_2D=>X"001000120010000B0004FFFCFFF5FFEFFFEDFFEFFFF3FFFA00020009000F0011",
		INIT_2E=>X"0007000E001200130010000A0002FFFAFFF2FFEEFFECFFEFFFF4FFFC0004000B",
		INIT_2F=>X"FFF800000009001000140013000F00080000FFF7FFF0FFECFFECFFEFFFF6FFFE",
		INIT_30=>X"FFEBFFF1FFFA0003000C001200150014000F0007FFFDFFF4FFEEFFEBFFEBFFF0",
		INIT_31=>X"FFE9FFE8FFEBFFF2FFFC0006000F001500160014000D0004FFFAFFF2FFEBFFE9",
		INIT_32=>X"FFF4FFECFFE7FFE7FFECFFF4FFFF00090012001700180014000C0002FFF7FFEF",
		INIT_33=>X"0008FFFCFFF0FFE8FFE5FFE6FFECFFF60002000D0015001900190013000AFFFF",
		INIT_34=>X"001A00110005FFF8FFECFFE5FFE2FFE6FFEEFFF9000500110018001B00190012",
		INIT_35=>X"001F0020001A000F0001FFF4FFE8FFE1FFE0FFE5FFEFFFFC00090015001C001E",
		INIT_36=>X"0013001E002300220019000CFFFDFFEFFFE3FFDEFFDEFFE5FFF10000000E0019",
		INIT_37=>X"FFF80009001900240027002300190009FFF8FFE9FFDEFFDAFFDDFFE6FFF40004",
		INIT_38=>X"FFD9FFE9FFFC00100020002A002C002500170005FFF3FFE3FFD8FFD6FFDBFFE7",
		INIT_39=>X"FFCAFFCCFFD8FFEB00020018002800310030002600150000FFECFFDBFFD2FFD1",
		INIT_3A=>X"FFD7FFC6FFC0FFC6FFD7FFEF000900220033003A003600280012FFFAFFE3FFD2",
		INIT_3B=>X"0008FFE5FFC8FFB6FFB3FFBEFFD5FFF40014002F00400045003D0029000EFFF1",
		INIT_3C=>X"0052002BFFFDFFD2FFB1FFA0FFA1FFB4FFD5FFFC00230042005300540045002A",
		INIT_3D=>X"00A200920067002BFFEBFFB2FF8AFF7AFF84FFA4FFD40009003B005F006F006A",
		INIT_3E=>X"00E0011E012100EF0097002CFFC2FF6DFF3AFF2FFF4BFF86FFD3002300680094",
		INIT_3F=>X"08F808AE07DA06940500034A01A0002CFF0DFE58FE0FFE29FE92FF2AFFD3006D",
		INIT_40=>X"0007000700050001FFFCFFF9FFF8FFF9FFFE00030006000700060002FFFDFFF9",
		INIT_41=>X"FFFBFFF8FFF8FFFBFFFF00040007000700050000FFFBFFF8FFF8FFFAFFFE0003",
		INIT_42=>X"00010005000700070003FFFFFFFAFFF8FFF8FFFB00000005000700070004FFFF",
		INIT_43=>X"0002FFFDFFF9FFF7FFF9FFFD00020006000800060003FFFEFFFAFFF8FFF8FFFC",
		INIT_44=>X"FFFAFFFE00030007000700050001FFFCFFF9FFF7FFF9FFFE0002000600080006",
		INIT_45=>X"00070004FFFFFFFBFFF8FFF8FFFBFFFF00040007000700050000FFFBFFF8FFF8",
		INIT_46=>X"FFF7FFF8FFFC00010005000700070003FFFFFFFAFFF8FFF8FFFB000000050007",
		INIT_47=>X"0006000800060002FFFDFFF9FFF7FFF9FFFD00020006000800060003FFFEFFFA",
		INIT_48=>X"FFFBFFF8FFF7FFFAFFFE00030007000800050001FFFCFFF8FFF7FFF9FFFD0002",
		INIT_49=>X"000000050007000700040000FFFBFFF8FFF8FFFAFFFF00040007000700050000",
		INIT_4A=>X"0003FFFEFFF9FFF7FFF8FFFC00010005000800070004FFFFFFFAFFF7FFF8FFFB",
		INIT_4B=>X"FFF9FFFD00020006000800060002FFFDFFF9FFF7FFF9FFFD0002000600080007",
		INIT_4C=>X"000800050000FFFBFFF8FFF7FFFAFFFE00030007000800060001FFFCFFF8FFF7",
		INIT_4D=>X"FFF7FFF8FFFB000000050008000800040000FFFBFFF8FFF7FFFAFFFF00040007",
		INIT_4E=>X"0006000800070003FFFEFFF9FFF7FFF8FFFC00010005000800070004FFFFFFFA",
		INIT_4F=>X"FFFCFFF8FFF7FFF9FFFD00020007000800060002FFFDFFF9FFF7FFF8FFFC0002",
		INIT_50=>X"FFFF00040008000800050001FFFBFFF8FFF7FFF9FFFE00030007000800060001",
		INIT_51=>X"0004FFFFFFFAFFF7FFF7FFFB000000050008000800050000FFFBFFF7FFF7FFFA",
		INIT_52=>X"FFF8FFFC00020006000800070003FFFEFFF9FFF7FFF8FFFB0001000600080008",
		INIT_53=>X"000900060002FFFCFFF8FFF6FFF8FFFD00020007000800070002FFFDFFF8FFF7",
		INIT_54=>X"FFF7FFF7FFFAFFFF00040008000800060001FFFBFFF7FFF6FFF9FFFE00030007",
		INIT_55=>X"0006000900080004FFFFFFFAFFF7FFF7FFFA000000050008000800050000FFFA",
		INIT_56=>X"FFFDFFF8FFF6FFF7FFFC00020006000900080004FFFEFFF9FFF6FFF7FFFB0001",
		INIT_57=>X"FFFE00030008000900070002FFFCFFF8FFF6FFF8FFFD00020007000900070003",
		INIT_58=>X"00060000FFFAFFF6FFF6FFF9FFFF00040008000900060001FFFBFFF7FFF6FFF8",
		INIT_59=>X"FFF6FFFB00010006000900090005FFFFFFF9FFF6FFF6FFFA0000000500090009",
		INIT_5A=>X"000A00080003FFFDFFF8FFF5FFF7FFFB00020007000900080004FFFEFFF9FFF6",
		INIT_5B=>X"FFF6FFF5FFF8FFFD00040008000A00070002FFFCFFF7FFF5FFF7FFFC00030008",
		INIT_5C=>X"00060009000A00060000FFFAFFF6FFF5FFF9FFFE00050009000A00070001FFFB",
		INIT_5D=>X"FFFEFFF8FFF5FFF6FFFA00010007000A00090005FFFFFFF9FFF5FFF5FFF9FFFF",
		INIT_5E=>X"FFFC00030008000A00090003FFFDFFF7FFF5FFF6FFFB00020007000A00090004",
		INIT_5F=>X"00080001FFFBFFF6FFF4FFF7FFFD00040009000B00080002FFFCFFF6FFF4FFF7",
		INIT_60=>X"FFF4FFF9FFFF0006000A000B00070000FFF9FFF5FFF4FFF8FFFE0005000A000B",
		INIT_61=>X"000B000A0005FFFEFFF7FFF4FFF5FFFA00010007000B000A0006FFFFFFF8FFF4",
		INIT_62=>X"FFF5FFF3FFF6FFFC00030009000C000A0004FFFDFFF6FFF4FFF5FFFA00020008",
		INIT_63=>X"0005000B000C00080002FFFAFFF5FFF3FFF6FFFD0004000A000C00090003FFFB",
		INIT_64=>X"FFFFFFF8FFF3FFF3FFF8FFFF0007000C000C00080000FFF9FFF4FFF3FFF7FFFE",
		INIT_65=>X"FFFA00020009000D000B0006FFFEFFF7FFF3FFF3FFF900000008000C000C0007",
		INIT_66=>X"000A0003FFFBFFF4FFF2FFF4FFFB0003000A000D000B0005FFFCFFF5FFF2FFF4",
		INIT_67=>X"FFF1FFF6FFFE0006000C000E000A0002FFFAFFF3FFF1FFF5FFFC0005000B000D",
		INIT_68=>X"000E000E0008FFFFFFF7FFF1FFF1FFF7FFFF0008000D000E00090001FFF8FFF2",
		INIT_69=>X"FFF4FFF0FFF2FFF90002000A000F000D0007FFFEFFF5FFF1FFF2FFF800000009",
		INIT_6A=>X"0005000D0010000C0004FFFAFFF3FFF0FFF2FFFA0004000C000F000D0006FFFC",
		INIT_6B=>X"0001FFF7FFF0FFEFFFF4FFFD0007000E0010000C0003FFF9FFF1FFEFFFF3FFFB",
		INIT_6C=>X"FFF60000000B00100010000AFFFFFFF5FFEFFFEFFFF5FFFF0009000F0010000B",
		INIT_6D=>X"00100007FFFCFFF2FFEDFFEFFFF70002000C001100100008FFFEFFF4FFEEFFEF",
		INIT_6E=>X"FFECFFF0FFFA000600100013000F0005FFFAFFF0FFECFFF0FFF90004000E0012",
		INIT_6F=>X"00130014000D0002FFF5FFEDFFEBFFF1FFFC000800110013000E0004FFF8FFEF",
		INIT_70=>X"FFF1FFEAFFEBFFF40000000D00140014000C0000FFF3FFEBFFEBFFF2FFFE000B",
		INIT_71=>X"00050011001700140009FFFBFFEFFFE9FFEBFFF50003000F00160014000BFFFD",
		INIT_72=>X"0005FFF6FFEAFFE6FFECFFF900080014001800130007FFF8FFECFFE7FFEBFFF7",
		INIT_73=>X"FFEEFFFE000E0018001A00120003FFF3FFE8FFE5FFEDFFFB000B001600190013",
		INIT_74=>X"001B000FFFFDFFECFFE3FFE4FFEF00000011001B001B00100000FFF0FFE5FFE5",
		INIT_75=>X"FFDFFFE4FFF300070018001F001B000DFFFAFFE9FFE1FFE4FFF100040014001D",
		INIT_76=>X"001F0024001B0008FFF2FFE2FFDCFFE4FFF6000B001B0021001B000AFFF6FFE5",
		INIT_77=>X"FFE9FFD9FFD8FFE6FFFC001400230026001A0004FFEEFFDEFFDAFFE5FFF9000F",
		INIT_78=>X"0005001F002C00290017FFFCFFE3FFD5FFD7FFE7000000190028002800190001",
		INIT_79=>X"0012FFF1FFD6FFCBFFD3FFEC000B00250032002B0015FFF7FFDDFFD0FFD5FFE9",
		INIT_7A=>X"FFD0FFF3001A0036003D002E000EFFE9FFCEFFC5FFD2FFEF0012002D0037002D",
		INIT_7B=>X"004E00310003FFD5FFB8FFB6FFCFFFF9002400410045002F0009FFE0FFC4FFBE",
		INIT_7C=>X"FF94FF9FFFCD000B0042006000590032FFFAFFC6FFA9FFACFFCE00000031004E",
		INIT_7D=>X"0082009E007E0033FFDAFF93FF77FF8DFFCC001A005B007800680033FFEDFFB1",
		INIT_7E=>X"FF6DFEF0FEE0FF37FFCB006400CB00E200A60034FFB8FF5FFF45FF70FFCB0034",
		INIT_7F=>X"0C980BCE099F068403280034FE2CFD4DFD85FE82FFCB00EA018A018A01030034",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_10,
		DOPADOP=>dopadop_10,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_11: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF003FFC00FFC00FFC00F",
		INITP_01=>X"FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FF000FFC00FFC00FFC",
		INITP_02=>X"C00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FF000FFC00FFC00",
		INITP_03=>X"0FFC00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF003FF000FFC00FF",
		INITP_04=>X"FC00FFC00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF003FFC00FFC0",
		INITP_05=>X"00FFC00FFC00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF003FFC00F",
		INITP_06=>X"FFC00FFC00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FF000FFC",
		INITP_07=>X"000FFC00FFC00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FF000",
		INITP_08=>X"FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC",
		INITP_09=>X"C03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00",
		INITP_0A=>X"0FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03F",
		INITP_0B=>X"FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F0",
		INITP_0C=>X"C0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00",
		INITP_0D=>X"0FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03F",
		INITP_0E=>X"FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F0",
		INITP_0F=>X"00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03",
		INIT_00=>X"0007000700050001FFFCFFF9FFF8FFF9FFFE00030006000700060002FFFDFFF9",
		INIT_01=>X"FFFBFFF8FFF8FFFBFFFF00040007000700050000FFFBFFF8FFF8FFFAFFFE0003",
		INIT_02=>X"00010005000700070003FFFFFFFAFFF8FFF8FFFB00000005000700070004FFFF",
		INIT_03=>X"0002FFFDFFF9FFF7FFF9FFFD00020006000800060003FFFEFFFAFFF8FFF8FFFC",
		INIT_04=>X"FFFAFFFE00030007000700050001FFFCFFF9FFF7FFF9FFFE0002000600080006",
		INIT_05=>X"00070004FFFFFFFBFFF8FFF8FFFBFFFF00040007000700050000FFFBFFF8FFF8",
		INIT_06=>X"FFF7FFF8FFFC00010005000700070003FFFFFFFAFFF8FFF8FFFB000000050007",
		INIT_07=>X"0006000800060002FFFDFFF9FFF7FFF9FFFD00020006000800060003FFFEFFFA",
		INIT_08=>X"FFFBFFF8FFF7FFFAFFFE00030007000800050001FFFCFFF8FFF7FFF9FFFD0002",
		INIT_09=>X"000000050007000700040000FFFBFFF8FFF8FFFAFFFF00040007000700050000",
		INIT_0A=>X"0003FFFEFFF9FFF7FFF8FFFC00010005000800070004FFFFFFFAFFF7FFF8FFFB",
		INIT_0B=>X"FFF9FFFD00020006000800060002FFFDFFF9FFF7FFF9FFFD0002000600080007",
		INIT_0C=>X"000800050000FFFBFFF8FFF7FFFAFFFE00030007000800060001FFFCFFF8FFF7",
		INIT_0D=>X"FFF7FFF8FFFB000000050008000800040000FFFBFFF8FFF7FFFAFFFF00040007",
		INIT_0E=>X"0006000800070003FFFEFFF9FFF7FFF8FFFC00010005000800070004FFFFFFFA",
		INIT_0F=>X"FFFCFFF8FFF7FFF9FFFD00020007000800060002FFFDFFF9FFF7FFF8FFFC0002",
		INIT_10=>X"FFFF00040008000800050001FFFBFFF8FFF7FFF9FFFE00030007000800060001",
		INIT_11=>X"0004FFFFFFFAFFF7FFF7FFFB000000050008000800050000FFFBFFF7FFF7FFFA",
		INIT_12=>X"FFF8FFFC00020006000800070003FFFEFFF9FFF7FFF8FFFB0001000600080008",
		INIT_13=>X"000900060002FFFCFFF8FFF6FFF8FFFD00020007000800070002FFFDFFF8FFF7",
		INIT_14=>X"FFF7FFF7FFFAFFFF00040008000800060001FFFBFFF7FFF6FFF9FFFE00030007",
		INIT_15=>X"0006000900080004FFFFFFFAFFF7FFF7FFFA000000050008000800050000FFFA",
		INIT_16=>X"FFFDFFF8FFF6FFF7FFFC00020006000900080004FFFEFFF9FFF6FFF7FFFB0001",
		INIT_17=>X"FFFE00030008000900070002FFFCFFF8FFF6FFF8FFFD00020007000900070003",
		INIT_18=>X"00060000FFFAFFF6FFF6FFF9FFFF00040008000900060001FFFBFFF7FFF6FFF8",
		INIT_19=>X"FFF6FFFB00010006000900090005FFFFFFF9FFF6FFF6FFFA0000000500090009",
		INIT_1A=>X"000A00080003FFFDFFF8FFF5FFF7FFFB00020007000900080004FFFEFFF9FFF6",
		INIT_1B=>X"FFF6FFF5FFF8FFFD00040008000A00070002FFFCFFF7FFF5FFF7FFFC00030008",
		INIT_1C=>X"00060009000A00060000FFFAFFF6FFF5FFF9FFFE00050009000A00070001FFFB",
		INIT_1D=>X"FFFEFFF8FFF5FFF6FFFA00010007000A00090005FFFFFFF9FFF5FFF5FFF9FFFF",
		INIT_1E=>X"FFFC00030008000A00090003FFFDFFF7FFF5FFF6FFFB00020007000A00090004",
		INIT_1F=>X"00080001FFFBFFF6FFF4FFF7FFFD00040009000B00080002FFFCFFF6FFF4FFF7",
		INIT_20=>X"FFF4FFF9FFFF0006000A000B00070000FFF9FFF5FFF4FFF8FFFE0005000A000B",
		INIT_21=>X"000B000A0005FFFEFFF7FFF4FFF5FFFA00010007000B000A0006FFFFFFF8FFF4",
		INIT_22=>X"FFF5FFF3FFF6FFFC00030009000C000A0004FFFDFFF6FFF4FFF5FFFA00020008",
		INIT_23=>X"0005000B000C00080002FFFAFFF5FFF3FFF6FFFD0004000A000C00090003FFFB",
		INIT_24=>X"FFFFFFF8FFF3FFF3FFF8FFFF0007000C000C00080000FFF9FFF4FFF3FFF7FFFE",
		INIT_25=>X"FFFA00020009000D000B0006FFFEFFF7FFF3FFF3FFF900000008000C000C0007",
		INIT_26=>X"000A0003FFFBFFF4FFF2FFF4FFFB0003000A000D000B0005FFFCFFF5FFF2FFF4",
		INIT_27=>X"FFF1FFF6FFFE0006000C000E000A0002FFFAFFF3FFF1FFF5FFFC0005000B000D",
		INIT_28=>X"000E000E0008FFFFFFF7FFF1FFF1FFF7FFFF0008000D000E00090001FFF8FFF2",
		INIT_29=>X"FFF4FFF0FFF2FFF90002000A000F000D0007FFFEFFF5FFF1FFF2FFF800000009",
		INIT_2A=>X"0005000D0010000C0004FFFAFFF3FFF0FFF2FFFA0004000C000F000D0006FFFC",
		INIT_2B=>X"0001FFF7FFF0FFEFFFF4FFFD0007000E0010000C0003FFF9FFF1FFEFFFF3FFFB",
		INIT_2C=>X"FFF60000000B00100010000AFFFFFFF5FFEFFFEFFFF5FFFF0009000F0010000B",
		INIT_2D=>X"00100007FFFCFFF2FFEDFFEFFFF70002000C001100100008FFFEFFF4FFEEFFEF",
		INIT_2E=>X"FFECFFF0FFFA000600100013000F0005FFFAFFF0FFECFFF0FFF90004000E0012",
		INIT_2F=>X"00130014000D0002FFF5FFEDFFEBFFF1FFFC000800110013000E0004FFF8FFEF",
		INIT_30=>X"FFF1FFEAFFEBFFF40000000D00140014000C0000FFF3FFEBFFEBFFF2FFFE000B",
		INIT_31=>X"00050011001700140009FFFBFFEFFFE9FFEBFFF50003000F00160014000BFFFD",
		INIT_32=>X"0005FFF6FFEAFFE6FFECFFF900080014001800130007FFF8FFECFFE7FFEBFFF7",
		INIT_33=>X"FFEEFFFE000E0018001A00120003FFF3FFE8FFE5FFEDFFFB000B001600190013",
		INIT_34=>X"001B000FFFFDFFECFFE3FFE4FFEF00000011001B001B00100000FFF0FFE5FFE5",
		INIT_35=>X"FFDFFFE4FFF300070018001F001B000DFFFAFFE9FFE1FFE4FFF100040014001D",
		INIT_36=>X"001F0024001B0008FFF2FFE2FFDCFFE4FFF6000B001B0021001B000AFFF6FFE5",
		INIT_37=>X"FFE9FFD9FFD8FFE6FFFC001400230026001A0004FFEEFFDEFFDAFFE5FFF9000F",
		INIT_38=>X"0005001F002C00290017FFFCFFE3FFD5FFD7FFE7000000190028002800190001",
		INIT_39=>X"0012FFF1FFD6FFCBFFD3FFEC000B00250032002B0015FFF7FFDDFFD0FFD5FFE9",
		INIT_3A=>X"FFD0FFF3001A0036003D002E000EFFE9FFCEFFC5FFD2FFEF0012002D0037002D",
		INIT_3B=>X"004E00310003FFD5FFB8FFB6FFCFFFF9002400410045002F0009FFE0FFC4FFBE",
		INIT_3C=>X"FF94FF9FFFCD000B0042006000590032FFFAFFC6FFA9FFACFFCE00000031004E",
		INIT_3D=>X"0082009E007E0033FFDAFF93FF77FF8DFFCC001A005B007800680033FFEDFFB1",
		INIT_3E=>X"FF6DFEF0FEE0FF37FFCB006400CB00E200A60034FFB8FF5FFF45FF70FFCB0034",
		INIT_3F=>X"0C980BCE099F068403280034FE2CFD4DFD85FE82FFCB00EA018A018A01030034",
		INIT_40=>X"0002000700070002FFFBFFF8FFFA0000000600070003FFFDFFF8FFF9FFFE0005",
		INIT_41=>X"FFF9FFFE000500080005FFFEFFF9FFF8FFFD0003000700060000FFFAFFF8FFFB",
		INIT_42=>X"FFFAFFF8FFFB0002000700070002FFFBFFF8FFFA0000000600070003FFFDFFF8",
		INIT_43=>X"0003FFFDFFF8FFF9FFFE000500080005FFFEFFF9FFF8FFFD0003000700060000",
		INIT_44=>X"000700060000FFFAFFF7FFFB0002000700070002FFFBFFF8FFFA000000060007",
		INIT_45=>X"0000000600070003FFFDFFF8FFF9FFFE000500080005FFFEFFF9FFF8FFFC0003",
		INIT_46=>X"FFF8FFFC0003000700060000FFFAFFF7FFFB0002000700070002FFFBFFF7FFFA",
		INIT_47=>X"FFFBFFF7FFFA0000000600070003FFFDFFF8FFF9FFFE000500080005FFFEFFF9",
		INIT_48=>X"0005FFFEFFF9FFF8FFFC0003000700060000FFFAFFF7FFFB0002000700070002",
		INIT_49=>X"000700070002FFFBFFF7FFF90000000600080003FFFDFFF8FFF8FFFE00050008",
		INIT_4A=>X"FFFE000500080005FFFEFFF8FFF8FFFC0003000800060000FFFAFFF7FFFB0002",
		INIT_4B=>X"FFF7FFFB0002000700070002FFFBFFF7FFF90000000600080003FFFCFFF8FFF8",
		INIT_4C=>X"FFFCFFF8FFF8FFFE000500080005FFFEFFF8FFF8FFFC0003000800060000FFF9",
		INIT_4D=>X"00060000FFF9FFF7FFFB0002000700070002FFFBFFF7FFF90000000600080004",
		INIT_4E=>X"000600080004FFFCFFF7FFF8FFFE000500080005FFFEFFF8FFF7FFFC00030008",
		INIT_4F=>X"FFFC0003000800060000FFF9FFF7FFFB0002000700070002FFFBFFF7FFF90000",
		INIT_50=>X"FFF7FFF90000000600080004FFFCFFF7FFF8FFFE000500080005FFFEFFF8FFF7",
		INIT_51=>X"FFFEFFF8FFF7FFFC0004000800070000FFF9FFF7FFFA0002000700080002FFFB",
		INIT_52=>X"00080002FFFBFFF7FFF90000000700080004FFFCFFF7FFF8FFFE000500080005",
		INIT_53=>X"000500090005FFFEFFF8FFF7FFFC0004000800070000FFF9FFF7FFFA00020008",
		INIT_54=>X"FFFA0002000800080002FFFAFFF6FFF90000000700080004FFFCFFF7FFF8FFFE",
		INIT_55=>X"FFF7FFF7FFFE000500090006FFFEFFF8FFF7FFFC0004000800070000FFF9FFF6",
		INIT_56=>X"0000FFF9FFF6FFFA0002000800080002FFFAFFF6FFF90000000700090004FFFC",
		INIT_57=>X"00090004FFFCFFF6FFF7FFFE000600090006FFFEFFF7FFF6FFFC000400090007",
		INIT_58=>X"0004000900070000FFF9FFF6FFFA0002000800080002FFFAFFF6FFF800000007",
		INIT_59=>X"FFF80000000700090004FFFCFFF6FFF7FFFE000600090006FFFEFFF7FFF6FFFC",
		INIT_5A=>X"FFF7FFF6FFFC0004000900080000FFF8FFF5FFFA0002000800090002FFFAFFF6",
		INIT_5B=>X"0003FFFAFFF5FFF800000008000A0005FFFCFFF6FFF7FFFE0006000A0006FFFE",
		INIT_5C=>X"000A0007FFFEFFF7FFF5FFFB0004000A00080000FFF8FFF5FFF9000200090009",
		INIT_5D=>X"0002000900090003FFFAFFF5FFF800000008000A0005FFFCFFF6FFF6FFFE0006",
		INIT_5E=>X"FFF6FFFD0006000A0007FFFEFFF6FFF5FFFB0004000A00080000FFF8FFF5FFF9",
		INIT_5F=>X"FFF8FFF4FFF90002000A000A0003FFF9FFF4FFF700000008000A0005FFFCFFF5",
		INIT_60=>X"0005FFFCFFF5FFF5FFFD0007000B0007FFFEFFF6FFF5FFFB0005000B00090000",
		INIT_61=>X"000B00090000FFF7FFF4FFF90002000A000A0003FFF9FFF4FFF700000009000B",
		INIT_62=>X"00000009000B0006FFFBFFF4FFF5FFFD0007000C0008FFFEFFF5FFF4FFFB0005",
		INIT_63=>X"FFF3FFFA0005000C000A0001FFF7FFF3FFF80002000B000B0003FFF9FFF3FFF6",
		INIT_64=>X"FFF9FFF3FFF60000000A000C0006FFFBFFF3FFF4FFFD0007000C0008FFFEFFF5",
		INIT_65=>X"0009FFFEFFF4FFF3FFFA0005000C000A0001FFF6FFF2FFF80003000B000C0003",
		INIT_66=>X"000C000C0004FFF8FFF2FFF50000000A000D0006FFFBFFF3FFF4FFFD0008000D",
		INIT_67=>X"FFFD0008000E0009FFFEFFF4FFF2FFFA0006000D000B0001FFF6FFF2FFF70003",
		INIT_68=>X"FFF1FFF70003000D000D0004FFF8FFF1FFF50000000B000E0007FFFBFFF2FFF3",
		INIT_69=>X"FFFAFFF1FFF2FFFC0009000F000AFFFEFFF3FFF1FFF90006000E000C0001FFF5",
		INIT_6A=>X"000D0001FFF4FFEFFFF60003000E000E0004FFF7FFF0FFF40000000C000F0007",
		INIT_6B=>X"000D00100008FFFAFFF0FFF1FFFC000A0010000BFFFDFFF2FFF0FFF90007000F",
		INIT_6C=>X"FFF800070011000E0001FFF3FFEEFFF50004000F000F0005FFF6FFEFFFF30000",
		INIT_6D=>X"FFEDFFF10000000E00120009FFF9FFEEFFF0FFFC000B0012000CFFFDFFF1FFEE",
		INIT_6E=>X"FFFDFFEFFFEDFFF800080012000F0001FFF2FFECFFF40004001000110005FFF6",
		INIT_6F=>X"00130006FFF5FFEBFFF00000000F0014000AFFF9FFEDFFEEFFFB000C0013000D",
		INIT_70=>X"000D0016000EFFFDFFEDFFEBFFF70009001400110002FFF1FFEAFFF300040012",
		INIT_71=>X"FFF10005001400150007FFF3FFE9FFEE000000110016000BFFF8FFEAFFECFFFB",
		INIT_72=>X"FFE8FFE9FFFA000F00190010FFFDFFEBFFE8FFF5000A001700130002FFEFFFE8",
		INIT_73=>X"0002FFECFFE4FFEF0006001700180008FFF2FFE5FFEC000000130019000DFFF7",
		INIT_74=>X"001D000FFFF6FFE4FFE6FFF90011001C0013FFFCFFE8FFE4FFF4000C001A0016",
		INIT_75=>X"000E001F001A0003FFE9FFE0FFED0007001B001C0009FFEFFFE1FFE800000017",
		INIT_76=>X"FFE40000001B00230012FFF4FFDFFFE1FFF8001500220017FFFCFFE4FFDFFFF2",
		INIT_77=>X"FFDDFFD8FFEF0011002600200003FFE5FFD9FFE9000800210022000BFFECFFDB",
		INIT_78=>X"000EFFE7FFD2FFDD00000022002B0016FFF1FFD7FFDAFFF700190029001CFFFB",
		INIT_79=>X"00360024FFF9FFD4FFCDFFEA0015003100290005FFDDFFCFFFE2000A002A002B",
		INIT_7A=>X"000E0039003B0013FFDFFFC3FFD10000002D0039001DFFEDFFCBFFCEFFF40021",
		INIT_7B=>X"FFB8FFEE0030004D0034FFF7FFC2FFB9FFE1001E004400390007FFD1FFBDFFD8",
		INIT_7C=>X"FFB5FF95FFC100160058005B001EFFCEFFA3FFBA000000430055002BFFE4FFB2",
		INIT_7D=>X"0053FFCDFF71FF7CFFE100550089005BFFF1FF96FF88FFCD0032006F005D000B",
		INIT_7E=>X"013A00FD001FFF43FEFBFF69003300C800C90042FF98FF41FF720000008400A6",
		INIT_7F=>X"11A80F860A0D0380FE5FFC36FD00FF60018A02420166FFCCFE98FE7DFF630092",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_11,
		DOPADOP=>dopadop_11,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_12: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC",
		INITP_01=>X"C03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00",
		INITP_02=>X"0FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03F",
		INITP_03=>X"FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F0",
		INITP_04=>X"C0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00",
		INITP_05=>X"0FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03F",
		INITP_06=>X"FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F0",
		INITP_07=>X"00FF03FC03F00FC03FC0FF00FC03F00FF03FC03F00FC03FC0FF00FC03F00FF03",
		INITP_08=>X"03F0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3",
		INITP_09=>X"3F03C0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0F",
		INITP_0A=>X"FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC",
		INITP_0B=>X"C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0",
		INITP_0C=>X"0FC3F03C0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3F03",
		INITP_0D=>X"3C0FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F",
		INITP_0E=>X"F03C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F0FC0F0",
		INITP_0F=>X"03F0FC3F03C0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3",
		INIT_00=>X"0002000700070002FFFBFFF8FFFA0000000600070003FFFDFFF8FFF9FFFE0005",
		INIT_01=>X"FFF9FFFE000500080005FFFEFFF9FFF8FFFD0003000700060000FFFAFFF8FFFB",
		INIT_02=>X"FFFAFFF8FFFB0002000700070002FFFBFFF8FFFA0000000600070003FFFDFFF8",
		INIT_03=>X"0003FFFDFFF8FFF9FFFE000500080005FFFEFFF9FFF8FFFD0003000700060000",
		INIT_04=>X"000700060000FFFAFFF7FFFB0002000700070002FFFBFFF8FFFA000000060007",
		INIT_05=>X"0000000600070003FFFDFFF8FFF9FFFE000500080005FFFEFFF9FFF8FFFC0003",
		INIT_06=>X"FFF8FFFC0003000700060000FFFAFFF7FFFB0002000700070002FFFBFFF7FFFA",
		INIT_07=>X"FFFBFFF7FFFA0000000600070003FFFDFFF8FFF9FFFE000500080005FFFEFFF9",
		INIT_08=>X"0005FFFEFFF9FFF8FFFC0003000700060000FFFAFFF7FFFB0002000700070002",
		INIT_09=>X"000700070002FFFBFFF7FFF90000000600080003FFFDFFF8FFF8FFFE00050008",
		INIT_0A=>X"FFFE000500080005FFFEFFF8FFF8FFFC0003000800060000FFFAFFF7FFFB0002",
		INIT_0B=>X"FFF7FFFB0002000700070002FFFBFFF7FFF90000000600080003FFFCFFF8FFF8",
		INIT_0C=>X"FFFCFFF8FFF8FFFE000500080005FFFEFFF8FFF8FFFC0003000800060000FFF9",
		INIT_0D=>X"00060000FFF9FFF7FFFB0002000700070002FFFBFFF7FFF90000000600080004",
		INIT_0E=>X"000600080004FFFCFFF7FFF8FFFE000500080005FFFEFFF8FFF7FFFC00030008",
		INIT_0F=>X"FFFC0003000800060000FFF9FFF7FFFB0002000700070002FFFBFFF7FFF90000",
		INIT_10=>X"FFF7FFF90000000600080004FFFCFFF7FFF8FFFE000500080005FFFEFFF8FFF7",
		INIT_11=>X"FFFEFFF8FFF7FFFC0004000800070000FFF9FFF7FFFA0002000700080002FFFB",
		INIT_12=>X"00080002FFFBFFF7FFF90000000700080004FFFCFFF7FFF8FFFE000500080005",
		INIT_13=>X"000500090005FFFEFFF8FFF7FFFC0004000800070000FFF9FFF7FFFA00020008",
		INIT_14=>X"FFFA0002000800080002FFFAFFF6FFF90000000700080004FFFCFFF7FFF8FFFE",
		INIT_15=>X"FFF7FFF7FFFE000500090006FFFEFFF8FFF7FFFC0004000800070000FFF9FFF6",
		INIT_16=>X"0000FFF9FFF6FFFA0002000800080002FFFAFFF6FFF90000000700090004FFFC",
		INIT_17=>X"00090004FFFCFFF6FFF7FFFE000600090006FFFEFFF7FFF6FFFC000400090007",
		INIT_18=>X"0004000900070000FFF9FFF6FFFA0002000800080002FFFAFFF6FFF800000007",
		INIT_19=>X"FFF80000000700090004FFFCFFF6FFF7FFFE000600090006FFFEFFF7FFF6FFFC",
		INIT_1A=>X"FFF7FFF6FFFC0004000900080000FFF8FFF5FFFA0002000800090002FFFAFFF6",
		INIT_1B=>X"0003FFFAFFF5FFF800000008000A0005FFFCFFF6FFF7FFFE0006000A0006FFFE",
		INIT_1C=>X"000A0007FFFEFFF7FFF5FFFB0004000A00080000FFF8FFF5FFF9000200090009",
		INIT_1D=>X"0002000900090003FFFAFFF5FFF800000008000A0005FFFCFFF6FFF6FFFE0006",
		INIT_1E=>X"FFF6FFFD0006000A0007FFFEFFF6FFF5FFFB0004000A00080000FFF8FFF5FFF9",
		INIT_1F=>X"FFF8FFF4FFF90002000A000A0003FFF9FFF4FFF700000008000A0005FFFCFFF5",
		INIT_20=>X"0005FFFCFFF5FFF5FFFD0007000B0007FFFEFFF6FFF5FFFB0005000B00090000",
		INIT_21=>X"000B00090000FFF7FFF4FFF90002000A000A0003FFF9FFF4FFF700000009000B",
		INIT_22=>X"00000009000B0006FFFBFFF4FFF5FFFD0007000C0008FFFEFFF5FFF4FFFB0005",
		INIT_23=>X"FFF3FFFA0005000C000A0001FFF7FFF3FFF80002000B000B0003FFF9FFF3FFF6",
		INIT_24=>X"FFF9FFF3FFF60000000A000C0006FFFBFFF3FFF4FFFD0007000C0008FFFEFFF5",
		INIT_25=>X"0009FFFEFFF4FFF3FFFA0005000C000A0001FFF6FFF2FFF80003000B000C0003",
		INIT_26=>X"000C000C0004FFF8FFF2FFF50000000A000D0006FFFBFFF3FFF4FFFD0008000D",
		INIT_27=>X"FFFD0008000E0009FFFEFFF4FFF2FFFA0006000D000B0001FFF6FFF2FFF70003",
		INIT_28=>X"FFF1FFF70003000D000D0004FFF8FFF1FFF50000000B000E0007FFFBFFF2FFF3",
		INIT_29=>X"FFFAFFF1FFF2FFFC0009000F000AFFFEFFF3FFF1FFF90006000E000C0001FFF5",
		INIT_2A=>X"000D0001FFF4FFEFFFF60003000E000E0004FFF7FFF0FFF40000000C000F0007",
		INIT_2B=>X"000D00100008FFFAFFF0FFF1FFFC000A0010000BFFFDFFF2FFF0FFF90007000F",
		INIT_2C=>X"FFF800070011000E0001FFF3FFEEFFF50004000F000F0005FFF6FFEFFFF30000",
		INIT_2D=>X"FFEDFFF10000000E00120009FFF9FFEEFFF0FFFC000B0012000CFFFDFFF1FFEE",
		INIT_2E=>X"FFFDFFEFFFEDFFF800080012000F0001FFF2FFECFFF40004001000110005FFF6",
		INIT_2F=>X"00130006FFF5FFEBFFF00000000F0014000AFFF9FFEDFFEEFFFB000C0013000D",
		INIT_30=>X"000D0016000EFFFDFFEDFFEBFFF70009001400110002FFF1FFEAFFF300040012",
		INIT_31=>X"FFF10005001400150007FFF3FFE9FFEE000000110016000BFFF8FFEAFFECFFFB",
		INIT_32=>X"FFE8FFE9FFFA000F00190010FFFDFFEBFFE8FFF5000A001700130002FFEFFFE8",
		INIT_33=>X"0002FFECFFE4FFEF0006001700180008FFF2FFE5FFEC000000130019000DFFF7",
		INIT_34=>X"001D000FFFF6FFE4FFE6FFF90011001C0013FFFCFFE8FFE4FFF4000C001A0016",
		INIT_35=>X"000E001F001A0003FFE9FFE0FFED0007001B001C0009FFEFFFE1FFE800000017",
		INIT_36=>X"FFE40000001B00230012FFF4FFDFFFE1FFF8001500220017FFFCFFE4FFDFFFF2",
		INIT_37=>X"FFDDFFD8FFEF0011002600200003FFE5FFD9FFE9000800210022000BFFECFFDB",
		INIT_38=>X"000EFFE7FFD2FFDD00000022002B0016FFF1FFD7FFDAFFF700190029001CFFFB",
		INIT_39=>X"00360024FFF9FFD4FFCDFFEA0015003100290005FFDDFFCFFFE2000A002A002B",
		INIT_3A=>X"000E0039003B0013FFDFFFC3FFD10000002D0039001DFFEDFFCBFFCEFFF40021",
		INIT_3B=>X"FFB8FFEE0030004D0034FFF7FFC2FFB9FFE1001E004400390007FFD1FFBDFFD8",
		INIT_3C=>X"FFB5FF95FFC100160058005B001EFFCEFFA3FFBA000000430055002BFFE4FFB2",
		INIT_3D=>X"0053FFCDFF71FF7CFFE100550089005BFFF1FF96FF88FFCD0032006F005D000B",
		INIT_3E=>X"013A00FD001FFF43FEFBFF69003300C800C90042FF98FF41FF720000008400A6",
		INIT_3F=>X"11A80F860A0D0380FE5FFC36FD00FF60018A02420166FFCCFE98FE7DFF630092",
		INIT_40=>X"FFF9FFF9000200070003FFFAFFF8000000070004FFFBFFF8FFFE00070006FFFD",
		INIT_41=>X"FFFCFFF8FFFD00060006FFFEFFF8FFFC00050007FFFFFFF8FFFA000300070001",
		INIT_42=>X"0000FFF8FFFA000200080002FFF9FFF9000100070004FFFBFFF8FFFF00070005",
		INIT_43=>X"0005FFFBFFF8FFFE00060006FFFDFFF7FFFC00050007FFFFFFF8FFFB00040007",
		INIT_44=>X"00070000FFF8FFFA000300080002FFF9FFF9000100070003FFFAFFF800000007",
		INIT_45=>X"00070004FFFBFFF8FFFF00070005FFFCFFF7FFFD00060006FFFEFFF8FFFB0005",
		INIT_46=>X"00050007FFFFFFF8FFFA000400070001FFF8FFF9000200080003FFFAFFF80000",
		INIT_47=>X"000100080004FFFAFFF8FFFF00070005FFFCFFF7FFFE00060006FFFDFFF7FFFC",
		INIT_48=>X"FFFD00060007FFFEFFF8FFFB000400070000FFF8FFFA000300080002FFF9FFF9",
		INIT_49=>X"FFF9000200080003FFFAFFF8000000070004FFFBFFF7FFFE00070006FFFDFFF7",
		INIT_4A=>X"FFF7FFFD00060006FFFEFFF7FFFC000500070000FFF8FFFA000300080001FFF9",
		INIT_4B=>X"FFF8FFF9000200080002FFF9FFF8000100080004FFFAFFF8FFFF00070005FFFC",
		INIT_4C=>X"FFFBFFF7FFFE00070006FFFDFFF7FFFC00060007FFFFFFF7FFFB000400080001",
		INIT_4D=>X"0000FFF8FFFA000300080002FFF9FFF8000100080003FFFAFFF8000000070005",
		INIT_4E=>X"0004FFFBFFF7FFFF00070006FFFCFFF7FFFD00060007FFFEFFF7FFFB00050008",
		INIT_4F=>X"0008FFFFFFF7FFFA000400080001FFF8FFF9000200080003FFF9FFF800000008",
		INIT_50=>X"00080004FFFAFFF7FFFF00080005FFFCFFF7FFFD00070007FFFDFFF7FFFC0005",
		INIT_51=>X"00060007FFFEFFF7FFFB000500080000FFF8FFF9000300080002FFF9FFF80001",
		INIT_52=>X"000200080003FFF9FFF7000000080005FFFBFFF7FFFE00070006FFFDFFF7FFFC",
		INIT_53=>X"FFFD00070007FFFEFFF7FFFB000500080000FFF7FFFA000400080002FFF8FFF8",
		INIT_54=>X"FFF9000300090003FFF9FFF7000100080004FFFAFFF7FFFF00080006FFFCFFF6",
		INIT_55=>X"FFF6FFFE00070007FFFDFFF6FFFC00060008FFFFFFF7FFFA000400090001FFF7",
		INIT_56=>X"FFF7FFF9000400090002FFF8FFF8000200090004FFF9FFF7000000080006FFFB",
		INIT_57=>X"FFFAFFF6FFFE00080007FFFCFFF6FFFC00070008FFFEFFF6FFFA000500090000",
		INIT_58=>X"FFFFFFF6FFF9000400090001FFF7FFF8000200090003FFF9FFF7000000090005",
		INIT_59=>X"0005FFF9FFF6FFFF00090006FFFBFFF6FFFD00080008FFFDFFF6FFFB00060009",
		INIT_5A=>X"0009FFFEFFF6FFFA000500090001FFF7FFF80003000A0003FFF8FFF700010009",
		INIT_5B=>X"000A0004FFF8FFF6000000090006FFFAFFF5FFFE00080007FFFCFFF5FFFC0007",
		INIT_5C=>X"00080008FFFDFFF5FFFA000600090000FFF6FFF80004000A0002FFF7FFF70002",
		INIT_5D=>X"0003000A0003FFF7FFF60001000A0005FFF9FFF5FFFF00090007FFFBFFF5FFFC",
		INIT_5E=>X"FFFD00090008FFFCFFF5FFFB00070009FFFFFFF5FFF90005000A0001FFF6FFF7",
		INIT_5F=>X"FFF80004000B0003FFF7FFF60002000B0005FFF8FFF5FFFF000A0007FFFAFFF5",
		INIT_60=>X"FFF4FFFE000A0008FFFBFFF4FFFC0008000AFFFEFFF4FFF90006000A0000FFF5",
		INIT_61=>X"FFF4FFF80005000B0002FFF5FFF60003000B0004FFF7FFF50000000B0006FFF9",
		INIT_62=>X"FFF8FFF4FFFF000B0008FFFAFFF3FFFC0009000AFFFDFFF4FFFA0007000BFFFF",
		INIT_63=>X"FFFEFFF3FFF80007000C0001FFF4FFF60004000C0004FFF6FFF50002000C0006",
		INIT_64=>X"0005FFF7FFF40000000C0008FFF9FFF3FFFD000A0009FFFCFFF3FFFB0009000B",
		INIT_65=>X"000BFFFDFFF2FFF90008000C0000FFF3FFF70005000D0003FFF5FFF50003000C",
		INIT_66=>X"000D0005FFF5FFF30001000D0007FFF8FFF2FFFE000C0009FFFAFFF2FFFB000A",
		INIT_67=>X"000B000BFFFCFFF1FFF90009000DFFFFFFF2FFF70007000D0002FFF3FFF50004",
		INIT_68=>X"0006000E0004FFF4FFF30002000E0007FFF6FFF2FFFF000D0009FFF9FFF1FFFC",
		INIT_69=>X"FFFD000D000BFFFAFFF0FFFA000B000DFFFDFFF1FFF70008000E0001FFF2FFF5",
		INIT_6A=>X"FFF50007000F0003FFF2FFF30004000F0006FFF4FFF10001000F0009FFF7FFF0",
		INIT_6B=>X"FFEFFFFE000F000BFFF8FFEFFFFB000D000DFFFCFFEFFFF8000A000FFFFFFFF0",
		INIT_6C=>X"FFEEFFF5000900110002FFF0FFF2000600110005FFF2FFF0000200100009FFF5",
		INIT_6D=>X"FFF3FFEE00000011000BFFF6FFEDFFFC000F000EFFFAFFEDFFF8000C0010FFFE",
		INIT_6E=>X"FFFCFFECFFF5000C00120000FFEEFFF2000800130004FFF0FFF0000400120008",
		INIT_6F=>X"0008FFF0FFED00020013000BFFF4FFECFFFD0012000EFFF8FFEBFFF9000F0011",
		INIT_70=>X"0012FFFAFFEAFFF6000E0014FFFFFFEBFFF2000B00150003FFEDFFEF00060014",
		INIT_71=>X"00170007FFEDFFEB00040016000BFFF1FFEAFFFF0015000FFFF5FFE9FFFA0012",
		INIT_72=>X"00160013FFF7FFE6FFF600120015FFFCFFE8FFF2000E00170002FFEAFFEE0009",
		INIT_73=>X"000C001B0006FFE9FFEA0007001A000BFFEDFFE700010018000FFFF2FFE6FFFB",
		INIT_74=>X"FFFD001B0015FFF3FFE2FFF700170018FFFAFFE3FFF20012001A0000FFE5FFED",
		INIT_75=>X"FFEC0011001F0004FFE3FFE7000B001F000AFFE8FFE40004001D0010FFEDFFE3",
		INIT_76=>X"FFDD000000210017FFEEFFDDFFF8001D001BFFF6FFDDFFF20018001EFFFDFFE0",
		INIT_77=>X"FFD7FFEA001800260002FFDBFFE400100026000AFFE1FFE0000800240011FFE7",
		INIT_78=>X"FFDEFFD60004002C001AFFE6FFD4FFFA00260020FFF0FFD5FFF100200024FFF9",
		INIT_79=>X"FFF2FFCAFFE700230030FFFEFFCFFFDF001900310009FFD6FFD9000E002F0012",
		INIT_7A=>X"0014FFCDFFC9000B003D001FFFD9FFC6FFFD00360027FFE6FFC7FFF1002D002D",
		INIT_7B=>X"003FFFE5FFB0FFE200380043FFF7FFB8FFD6002900440007FFC2FFCE00190042",
		INIT_7C=>X"006B0018FFA9FFAC001A0062002AFFBEFFAA000400550036FFD2FFABFFF10047",
		INIT_7D=>X"00930071FFC2FF6BFFD5006F0074FFE5FF7FFFC1004F00720002FF94FFB40033",
		INIT_7E=>X"00AE012C002BFF10FF39005400ED0051FF5DFF47001A00BC0066FF95FF58FFF1",
		INIT_7F=>X"18B8131506ADFCC0FAF5FF2002DA0255FF4AFDBEFF25014D018CFFE5FE9BFF2D",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_12,
		DOPADOP=>dopadop_12,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_13: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"03F0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3",
		INITP_01=>X"3F03C0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0F",
		INITP_02=>X"FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC",
		INITP_03=>X"C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0",
		INITP_04=>X"0FC3F03C0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3F03",
		INITP_05=>X"3C0FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F",
		INITP_06=>X"F03C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0F03F0FC3F0FC0F0",
		INITP_07=>X"03F0FC3F03C0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3",
		INITP_08=>X"F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F",
		INITP_09=>X"C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0",
		INITP_0A=>X"3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3",
		INITP_0B=>X"F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C",
		INITP_0C=>X"CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0",
		INITP_0D=>X"3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3",
		INITP_0E=>X"F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C",
		INITP_0F=>X"0F0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0",
		INIT_00=>X"FFF9FFF9000200070003FFFAFFF8000000070004FFFBFFF8FFFE00070006FFFD",
		INIT_01=>X"FFFCFFF8FFFD00060006FFFEFFF8FFFC00050007FFFFFFF8FFFA000300070001",
		INIT_02=>X"0000FFF8FFFA000200080002FFF9FFF9000100070004FFFBFFF8FFFF00070005",
		INIT_03=>X"0005FFFBFFF8FFFE00060006FFFDFFF7FFFC00050007FFFFFFF8FFFB00040007",
		INIT_04=>X"00070000FFF8FFFA000300080002FFF9FFF9000100070003FFFAFFF800000007",
		INIT_05=>X"00070004FFFBFFF8FFFF00070005FFFCFFF7FFFD00060006FFFEFFF8FFFB0005",
		INIT_06=>X"00050007FFFFFFF8FFFA000400070001FFF8FFF9000200080003FFFAFFF80000",
		INIT_07=>X"000100080004FFFAFFF8FFFF00070005FFFCFFF7FFFE00060006FFFDFFF7FFFC",
		INIT_08=>X"FFFD00060007FFFEFFF8FFFB000400070000FFF8FFFA000300080002FFF9FFF9",
		INIT_09=>X"FFF9000200080003FFFAFFF8000000070004FFFBFFF7FFFE00070006FFFDFFF7",
		INIT_0A=>X"FFF7FFFD00060006FFFEFFF7FFFC000500070000FFF8FFFA000300080001FFF9",
		INIT_0B=>X"FFF8FFF9000200080002FFF9FFF8000100080004FFFAFFF8FFFF00070005FFFC",
		INIT_0C=>X"FFFBFFF7FFFE00070006FFFDFFF7FFFC00060007FFFFFFF7FFFB000400080001",
		INIT_0D=>X"0000FFF8FFFA000300080002FFF9FFF8000100080003FFFAFFF8000000070005",
		INIT_0E=>X"0004FFFBFFF7FFFF00070006FFFCFFF7FFFD00060007FFFEFFF7FFFB00050008",
		INIT_0F=>X"0008FFFFFFF7FFFA000400080001FFF8FFF9000200080003FFF9FFF800000008",
		INIT_10=>X"00080004FFFAFFF7FFFF00080005FFFCFFF7FFFD00070007FFFDFFF7FFFC0005",
		INIT_11=>X"00060007FFFEFFF7FFFB000500080000FFF8FFF9000300080002FFF9FFF80001",
		INIT_12=>X"000200080003FFF9FFF7000000080005FFFBFFF7FFFE00070006FFFDFFF7FFFC",
		INIT_13=>X"FFFD00070007FFFEFFF7FFFB000500080000FFF7FFFA000400080002FFF8FFF8",
		INIT_14=>X"FFF9000300090003FFF9FFF7000100080004FFFAFFF7FFFF00080006FFFCFFF6",
		INIT_15=>X"FFF6FFFE00070007FFFDFFF6FFFC00060008FFFFFFF7FFFA000400090001FFF7",
		INIT_16=>X"FFF7FFF9000400090002FFF8FFF8000200090004FFF9FFF7000000080006FFFB",
		INIT_17=>X"FFFAFFF6FFFE00080007FFFCFFF6FFFC00070008FFFEFFF6FFFA000500090000",
		INIT_18=>X"FFFFFFF6FFF9000400090001FFF7FFF8000200090003FFF9FFF7000000090005",
		INIT_19=>X"0005FFF9FFF6FFFF00090006FFFBFFF6FFFD00080008FFFDFFF6FFFB00060009",
		INIT_1A=>X"0009FFFEFFF6FFFA000500090001FFF7FFF80003000A0003FFF8FFF700010009",
		INIT_1B=>X"000A0004FFF8FFF6000000090006FFFAFFF5FFFE00080007FFFCFFF5FFFC0007",
		INIT_1C=>X"00080008FFFDFFF5FFFA000600090000FFF6FFF80004000A0002FFF7FFF70002",
		INIT_1D=>X"0003000A0003FFF7FFF60001000A0005FFF9FFF5FFFF00090007FFFBFFF5FFFC",
		INIT_1E=>X"FFFD00090008FFFCFFF5FFFB00070009FFFFFFF5FFF90005000A0001FFF6FFF7",
		INIT_1F=>X"FFF80004000B0003FFF7FFF60002000B0005FFF8FFF5FFFF000A0007FFFAFFF5",
		INIT_20=>X"FFF4FFFE000A0008FFFBFFF4FFFC0008000AFFFEFFF4FFF90006000A0000FFF5",
		INIT_21=>X"FFF4FFF80005000B0002FFF5FFF60003000B0004FFF7FFF50000000B0006FFF9",
		INIT_22=>X"FFF8FFF4FFFF000B0008FFFAFFF3FFFC0009000AFFFDFFF4FFFA0007000BFFFF",
		INIT_23=>X"FFFEFFF3FFF80007000C0001FFF4FFF60004000C0004FFF6FFF50002000C0006",
		INIT_24=>X"0005FFF7FFF40000000C0008FFF9FFF3FFFD000A0009FFFCFFF3FFFB0009000B",
		INIT_25=>X"000BFFFDFFF2FFF90008000C0000FFF3FFF70005000D0003FFF5FFF50003000C",
		INIT_26=>X"000D0005FFF5FFF30001000D0007FFF8FFF2FFFE000C0009FFFAFFF2FFFB000A",
		INIT_27=>X"000B000BFFFCFFF1FFF90009000DFFFFFFF2FFF70007000D0002FFF3FFF50004",
		INIT_28=>X"0006000E0004FFF4FFF30002000E0007FFF6FFF2FFFF000D0009FFF9FFF1FFFC",
		INIT_29=>X"FFFD000D000BFFFAFFF0FFFA000B000DFFFDFFF1FFF70008000E0001FFF2FFF5",
		INIT_2A=>X"FFF50007000F0003FFF2FFF30004000F0006FFF4FFF10001000F0009FFF7FFF0",
		INIT_2B=>X"FFEFFFFE000F000BFFF8FFEFFFFB000D000DFFFCFFEFFFF8000A000FFFFFFFF0",
		INIT_2C=>X"FFEEFFF5000900110002FFF0FFF2000600110005FFF2FFF0000200100009FFF5",
		INIT_2D=>X"FFF3FFEE00000011000BFFF6FFEDFFFC000F000EFFFAFFEDFFF8000C0010FFFE",
		INIT_2E=>X"FFFCFFECFFF5000C00120000FFEEFFF2000800130004FFF0FFF0000400120008",
		INIT_2F=>X"0008FFF0FFED00020013000BFFF4FFECFFFD0012000EFFF8FFEBFFF9000F0011",
		INIT_30=>X"0012FFFAFFEAFFF6000E0014FFFFFFEBFFF2000B00150003FFEDFFEF00060014",
		INIT_31=>X"00170007FFEDFFEB00040016000BFFF1FFEAFFFF0015000FFFF5FFE9FFFA0012",
		INIT_32=>X"00160013FFF7FFE6FFF600120015FFFCFFE8FFF2000E00170002FFEAFFEE0009",
		INIT_33=>X"000C001B0006FFE9FFEA0007001A000BFFEDFFE700010018000FFFF2FFE6FFFB",
		INIT_34=>X"FFFD001B0015FFF3FFE2FFF700170018FFFAFFE3FFF20012001A0000FFE5FFED",
		INIT_35=>X"FFEC0011001F0004FFE3FFE7000B001F000AFFE8FFE40004001D0010FFEDFFE3",
		INIT_36=>X"FFDD000000210017FFEEFFDDFFF8001D001BFFF6FFDDFFF20018001EFFFDFFE0",
		INIT_37=>X"FFD7FFEA001800260002FFDBFFE400100026000AFFE1FFE0000800240011FFE7",
		INIT_38=>X"FFDEFFD60004002C001AFFE6FFD4FFFA00260020FFF0FFD5FFF100200024FFF9",
		INIT_39=>X"FFF2FFCAFFE700230030FFFEFFCFFFDF001900310009FFD6FFD9000E002F0012",
		INIT_3A=>X"0014FFCDFFC9000B003D001FFFD9FFC6FFFD00360027FFE6FFC7FFF1002D002D",
		INIT_3B=>X"003FFFE5FFB0FFE200380043FFF7FFB8FFD6002900440007FFC2FFCE00190042",
		INIT_3C=>X"006B0018FFA9FFAC001A0062002AFFBEFFAA000400550036FFD2FFABFFF10047",
		INIT_3D=>X"00930071FFC2FF6BFFD5006F0074FFE5FF7FFFC1004F00720002FF94FFB40033",
		INIT_3E=>X"00AE012C002BFF10FF39005400ED0051FF5DFF47001A00BC0066FF95FF58FFF1",
		INIT_3F=>X"18B8131506ADFCC0FAF5FF2002DA0255FF4AFDBEFF25014D018CFFE5FE9BFF2D",
		INIT_40=>X"FFFC00070002FFF800000007FFFDFFF800040006FFFAFFFB00060003FFF8FFFE",
		INIT_41=>X"FFFBFFF900050004FFF9FFFD00070000FFF700010007FFFCFFF900040005FFF9",
		INIT_42=>X"0008FFFEFFF800030006FFFAFFFA00060003FFF8FFFE0007FFFFFFF800020007",
		INIT_43=>X"FFFC00070001FFF800000007FFFDFFF800040006FFFAFFFB00070002FFF8FFFF",
		INIT_44=>X"FFFBFFF900050004FFF8FFFD00070000FFF700010007FFFCFFF900050005FFF9",
		INIT_45=>X"0008FFFEFFF800030006FFFAFFFA00060003FFF8FFFE0008FFFFFFF800020007",
		INIT_46=>X"FFFC00070001FFF700000007FFFDFFF800040006FFF9FFFB00070002FFF8FFFF",
		INIT_47=>X"FFFBFFF900060004FFF8FFFD00070000FFF700010007FFFCFFF900050005FFF9",
		INIT_48=>X"0008FFFEFFF800030006FFFAFFFA00060003FFF8FFFE0008FFFFFFF700020007",
		INIT_49=>X"FFFC00070001FFF700000008FFFDFFF800040006FFF9FFFB00070002FFF7FFFF",
		INIT_4A=>X"FFFBFFF900060004FFF8FFFD00080000FFF700010007FFFCFFF900050005FFF9",
		INIT_4B=>X"0008FFFEFFF800030006FFFAFFFA00070003FFF8FFFE0008FFFFFFF700020007",
		INIT_4C=>X"FFFC00080001FFF700000008FFFDFFF800040006FFF9FFFB00070002FFF7FFFF",
		INIT_4D=>X"FFFAFFF900060004FFF8FFFD00080000FFF700020007FFFBFFF900050005FFF8",
		INIT_4E=>X"0008FFFDFFF800040006FFFAFFFA00070003FFF7FFFE0008FFFFFFF700030007",
		INIT_4F=>X"FFFC00080001FFF700010008FFFCFFF800050006FFF9FFFB00070002FFF7FFFF",
		INIT_50=>X"FFFAFFF900060004FFF7FFFD0008FFFFFFF700020008FFFBFFF900060005FFF8",
		INIT_51=>X"0008FFFDFFF700040006FFF9FFFA00070003FFF7FFFE0008FFFEFFF700030007",
		INIT_52=>X"FFFC00080000FFF700010008FFFCFFF800050006FFF8FFFB00080002FFF70000",
		INIT_53=>X"FFFAFFF900070004FFF7FFFD0008FFFFFFF700020008FFFBFFF900060005FFF8",
		INIT_54=>X"0009FFFDFFF700040007FFF9FFFA00080003FFF7FFFF0009FFFEFFF700030007",
		INIT_55=>X"FFFC00090000FFF600010008FFFCFFF800050006FFF8FFFB00080002FFF60000",
		INIT_56=>X"FFF9FFF900070004FFF7FFFE0009FFFFFFF600020008FFFAFFF800060005FFF7",
		INIT_57=>X"0009FFFCFFF700050007FFF8FFFA00080003FFF6FFFF0009FFFEFFF600040007",
		INIT_58=>X"FFFC00090000FFF600010009FFFBFFF700060006FFF7FFFB00090001FFF60000",
		INIT_59=>X"FFF9FFF900080004FFF6FFFE0009FFFFFFF600030008FFFAFFF800070005FFF7",
		INIT_5A=>X"0009FFFCFFF700050007FFF8FFFA00090003FFF6FFFF0009FFFDFFF600040008",
		INIT_5B=>X"FFFC000A0000FFF500020009FFFBFFF700060006FFF7FFFB00090001FFF50000",
		INIT_5C=>X"FFF8FFF900080004FFF5FFFE000AFFFEFFF500030009FFF9FFF800080005FFF6",
		INIT_5D=>X"000AFFFCFFF600060007FFF7FFFA00090002FFF5FFFF000AFFFDFFF600050008",
		INIT_5E=>X"FFFD000A0000FFF50002000AFFFAFFF700070006FFF6FFFB000A0001FFF50001",
		INIT_5F=>X"FFF8FFF900090004FFF5FFFE000BFFFEFFF500040009FFF9FFF800080005FFF5",
		INIT_60=>X"000BFFFBFFF600070008FFF6FFFA000A0002FFF40000000BFFFDFFF500050008",
		INIT_61=>X"FFFD000BFFFFFFF40003000AFFF9FFF600080007FFF5FFFB000B0001FFF40001",
		INIT_62=>X"FFF7FFF8000A0004FFF4FFFE000CFFFEFFF40004000AFFF8FFF700090005FFF4",
		INIT_63=>X"000CFFFAFFF500070008FFF5FFFA000B0002FFF30000000CFFFCFFF400060009",
		INIT_64=>X"FFFD000CFFFFFFF30003000BFFF9FFF600090007FFF4FFFB000C0001FFF30002",
		INIT_65=>X"FFF6FFF8000B0004FFF2FFFE000DFFFDFFF30005000BFFF7FFF7000A0006FFF3",
		INIT_66=>X"000DFFF9FFF400090009FFF4FFF9000C0002FFF20000000DFFFBFFF30007000A",
		INIT_67=>X"FFFD000EFFFFFFF10004000CFFF8FFF5000A0007FFF3FFFB000D0001FFF20002",
		INIT_68=>X"FFF4FFF7000D0004FFF1FFFF000EFFFDFFF20006000CFFF6FFF6000C0006FFF2",
		INIT_69=>X"000EFFF8FFF3000A0009FFF3FFF9000E0002FFF00001000EFFFBFFF20008000B",
		INIT_6A=>X"FFFD0010FFFEFFF00005000EFFF6FFF4000C0008FFF1FFFB000F0000FFF00003",
		INIT_6B=>X"FFF2FFF7000F0004FFEFFFFF0010FFFCFFF00007000DFFF4FFF5000D0006FFF0",
		INIT_6C=>X"0010FFF7FFF1000C000BFFF1FFF800100002FFEE00010010FFF9FFF00009000C",
		INIT_6D=>X"FFFD0012FFFDFFEE00060010FFF5FFF2000E0009FFEFFFFA00110000FFEE0004",
		INIT_6E=>X"FFF0FFF600120005FFECFFFF0013FFFBFFEE0009000FFFF2FFF400100007FFED",
		INIT_6F=>X"0013FFF5FFEF000E000CFFEEFFF800130002FFEB00020013FFF8FFEE000B000E",
		INIT_70=>X"FFFD0016FFFCFFEA00080012FFF2FFF00011000AFFECFFFA0015FFFFFFEB0005",
		INIT_71=>X"FFECFFF400150005FFE800000016FFF9FFEA000B0011FFEFFFF200130008FFEA",
		INIT_72=>X"0017FFF2FFEC0012000EFFEAFFF600170002FFE700030017FFF6FFEB000E0010",
		INIT_73=>X"FFFD001BFFFBFFE6000B0016FFEFFFED0015000CFFE7FFF90019FFFFFFE60007",
		INIT_74=>X"FFE7FFF2001B0006FFE20001001CFFF7FFE5000F0015FFEBFFEF00180009FFE5",
		INIT_75=>X"001DFFEEFFE700170012FFE3FFF5001E0002FFE00005001DFFF3FFE600130014",
		INIT_76=>X"FFFD0024FFF9FFDE000F001DFFE9FFE8001C000FFFDFFFF80021FFFEFFDF000A",
		INIT_77=>X"FFDDFFED00260007FFD800020026FFF3FFDD0015001CFFE3FFEA0021000CFFDB",
		INIT_78=>X"0029FFE5FFDD00220018FFD7FFF1002B0002FFD400080028FFEDFFDD001B001B",
		INIT_79=>X"FFFD0035FFF4FFCE0017002AFFDDFFDE002A0015FFD1FFF60030FFFCFFD1000F",
		INIT_7A=>X"FFC8FFE4003C000AFFC10005003BFFEBFFCB0021002AFFD4FFE100320010FFC9",
		INIT_7B=>X"0047FFD1FFC6003C0028FFBBFFEA00480002FFB8000F0041FFDFFFC8002D002A",
		INIT_7C=>X"FFFD0069FFE7FFA0002F004FFFBDFFC4004F0025FFA9FFF10057FFF7FFAD001D",
		INIT_7D=>X"FF74FFC100930016FF6F000F0085FFCFFF8D004B0059FFA1FFC2006A001FFF92",
		INIT_7E=>X"011BFF47FF3100D80084FF1BFFC000E00002FF30003100B3FFA5FF6F00790068",
		INIT_7F=>X"22A81432FD5FF9B80289033DFD9BFE38023300E0FE08FFBF01B2FFCEFE970082",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_13,
		DOPADOP=>dopadop_13,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_14: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F",
		INITP_01=>X"C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0",
		INITP_02=>X"3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3",
		INITP_03=>X"F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C",
		INITP_04=>X"CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0",
		INITP_05=>X"3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3CF0F0F0C3C3C30F0F0F3C3C3",
		INITP_06=>X"F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C",
		INITP_07=>X"0F0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0F0C3C3C3CF0F0F3C3C3C30F0",
		INITP_08=>X"C33CCF30CF30CF30CF33CC33CC33CC33CCF30CF30CF30CF30CC33CC33CC33CC3",
		INITP_09=>X"3CC33CC330CF30CF30CF30CC33CC33CC33CC330CF30CF30CF30CF33CC33CC33C",
		INITP_0A=>X"C33CC33CC33CCF30CF30CF30CF33CC33CC33CC33CCF30CF30CF30CF33CC33CC3",
		INITP_0B=>X"3CC33CC33CC33CC330CF30CF30CF30CC33CC33CC33CC330CF30CF30CF30CC33C",
		INITP_0C=>X"F30CC33CC33CC33CC330CF30CF30CF30CF33CC33CC33CC33CCF30CF30CF30CF3",
		INITP_0D=>X"0CF30CF33CC33CC33CC33CCF30CF30CF30CF30CC33CC33CC33CC330CF30CF30C",
		INITP_0E=>X"F30CF30CF30CC33CC33CC33CC330CF30CF30CF30CC33CC33CC33CC33CCF30CF3",
		INITP_0F=>X"0CF30CF30CF30CF33CC33CC33CC33CCF30CF30CF30CF33CC33CC33CC33CC330C",
		INIT_00=>X"FFFC00070002FFF800000007FFFDFFF800040006FFFAFFFB00060003FFF8FFFE",
		INIT_01=>X"FFFBFFF900050004FFF9FFFD00070000FFF700010007FFFCFFF900040005FFF9",
		INIT_02=>X"0008FFFEFFF800030006FFFAFFFA00060003FFF8FFFE0007FFFFFFF800020007",
		INIT_03=>X"FFFC00070001FFF800000007FFFDFFF800040006FFFAFFFB00070002FFF8FFFF",
		INIT_04=>X"FFFBFFF900050004FFF8FFFD00070000FFF700010007FFFCFFF900050005FFF9",
		INIT_05=>X"0008FFFEFFF800030006FFFAFFFA00060003FFF8FFFE0008FFFFFFF800020007",
		INIT_06=>X"FFFC00070001FFF700000007FFFDFFF800040006FFF9FFFB00070002FFF8FFFF",
		INIT_07=>X"FFFBFFF900060004FFF8FFFD00070000FFF700010007FFFCFFF900050005FFF9",
		INIT_08=>X"0008FFFEFFF800030006FFFAFFFA00060003FFF8FFFE0008FFFFFFF700020007",
		INIT_09=>X"FFFC00070001FFF700000008FFFDFFF800040006FFF9FFFB00070002FFF7FFFF",
		INIT_0A=>X"FFFBFFF900060004FFF8FFFD00080000FFF700010007FFFCFFF900050005FFF9",
		INIT_0B=>X"0008FFFEFFF800030006FFFAFFFA00070003FFF8FFFE0008FFFFFFF700020007",
		INIT_0C=>X"FFFC00080001FFF700000008FFFDFFF800040006FFF9FFFB00070002FFF7FFFF",
		INIT_0D=>X"FFFAFFF900060004FFF8FFFD00080000FFF700020007FFFBFFF900050005FFF8",
		INIT_0E=>X"0008FFFDFFF800040006FFFAFFFA00070003FFF7FFFE0008FFFFFFF700030007",
		INIT_0F=>X"FFFC00080001FFF700010008FFFCFFF800050006FFF9FFFB00070002FFF7FFFF",
		INIT_10=>X"FFFAFFF900060004FFF7FFFD0008FFFFFFF700020008FFFBFFF900060005FFF8",
		INIT_11=>X"0008FFFDFFF700040006FFF9FFFA00070003FFF7FFFE0008FFFEFFF700030007",
		INIT_12=>X"FFFC00080000FFF700010008FFFCFFF800050006FFF8FFFB00080002FFF70000",
		INIT_13=>X"FFFAFFF900070004FFF7FFFD0008FFFFFFF700020008FFFBFFF900060005FFF8",
		INIT_14=>X"0009FFFDFFF700040007FFF9FFFA00080003FFF7FFFF0009FFFEFFF700030007",
		INIT_15=>X"FFFC00090000FFF600010008FFFCFFF800050006FFF8FFFB00080002FFF60000",
		INIT_16=>X"FFF9FFF900070004FFF7FFFE0009FFFFFFF600020008FFFAFFF800060005FFF7",
		INIT_17=>X"0009FFFCFFF700050007FFF8FFFA00080003FFF6FFFF0009FFFEFFF600040007",
		INIT_18=>X"FFFC00090000FFF600010009FFFBFFF700060006FFF7FFFB00090001FFF60000",
		INIT_19=>X"FFF9FFF900080004FFF6FFFE0009FFFFFFF600030008FFFAFFF800070005FFF7",
		INIT_1A=>X"0009FFFCFFF700050007FFF8FFFA00090003FFF6FFFF0009FFFDFFF600040008",
		INIT_1B=>X"FFFC000A0000FFF500020009FFFBFFF700060006FFF7FFFB00090001FFF50000",
		INIT_1C=>X"FFF8FFF900080004FFF5FFFE000AFFFEFFF500030009FFF9FFF800080005FFF6",
		INIT_1D=>X"000AFFFCFFF600060007FFF7FFFA00090002FFF5FFFF000AFFFDFFF600050008",
		INIT_1E=>X"FFFD000A0000FFF50002000AFFFAFFF700070006FFF6FFFB000A0001FFF50001",
		INIT_1F=>X"FFF8FFF900090004FFF5FFFE000BFFFEFFF500040009FFF9FFF800080005FFF5",
		INIT_20=>X"000BFFFBFFF600070008FFF6FFFA000A0002FFF40000000BFFFDFFF500050008",
		INIT_21=>X"FFFD000BFFFFFFF40003000AFFF9FFF600080007FFF5FFFB000B0001FFF40001",
		INIT_22=>X"FFF7FFF8000A0004FFF4FFFE000CFFFEFFF40004000AFFF8FFF700090005FFF4",
		INIT_23=>X"000CFFFAFFF500070008FFF5FFFA000B0002FFF30000000CFFFCFFF400060009",
		INIT_24=>X"FFFD000CFFFFFFF30003000BFFF9FFF600090007FFF4FFFB000C0001FFF30002",
		INIT_25=>X"FFF6FFF8000B0004FFF2FFFE000DFFFDFFF30005000BFFF7FFF7000A0006FFF3",
		INIT_26=>X"000DFFF9FFF400090009FFF4FFF9000C0002FFF20000000DFFFBFFF30007000A",
		INIT_27=>X"FFFD000EFFFFFFF10004000CFFF8FFF5000A0007FFF3FFFB000D0001FFF20002",
		INIT_28=>X"FFF4FFF7000D0004FFF1FFFF000EFFFDFFF20006000CFFF6FFF6000C0006FFF2",
		INIT_29=>X"000EFFF8FFF3000A0009FFF3FFF9000E0002FFF00001000EFFFBFFF20008000B",
		INIT_2A=>X"FFFD0010FFFEFFF00005000EFFF6FFF4000C0008FFF1FFFB000F0000FFF00003",
		INIT_2B=>X"FFF2FFF7000F0004FFEFFFFF0010FFFCFFF00007000DFFF4FFF5000D0006FFF0",
		INIT_2C=>X"0010FFF7FFF1000C000BFFF1FFF800100002FFEE00010010FFF9FFF00009000C",
		INIT_2D=>X"FFFD0012FFFDFFEE00060010FFF5FFF2000E0009FFEFFFFA00110000FFEE0004",
		INIT_2E=>X"FFF0FFF600120005FFECFFFF0013FFFBFFEE0009000FFFF2FFF400100007FFED",
		INIT_2F=>X"0013FFF5FFEF000E000CFFEEFFF800130002FFEB00020013FFF8FFEE000B000E",
		INIT_30=>X"FFFD0016FFFCFFEA00080012FFF2FFF00011000AFFECFFFA0015FFFFFFEB0005",
		INIT_31=>X"FFECFFF400150005FFE800000016FFF9FFEA000B0011FFEFFFF200130008FFEA",
		INIT_32=>X"0017FFF2FFEC0012000EFFEAFFF600170002FFE700030017FFF6FFEB000E0010",
		INIT_33=>X"FFFD001BFFFBFFE6000B0016FFEFFFED0015000CFFE7FFF90019FFFFFFE60007",
		INIT_34=>X"FFE7FFF2001B0006FFE20001001CFFF7FFE5000F0015FFEBFFEF00180009FFE5",
		INIT_35=>X"001DFFEEFFE700170012FFE3FFF5001E0002FFE00005001DFFF3FFE600130014",
		INIT_36=>X"FFFD0024FFF9FFDE000F001DFFE9FFE8001C000FFFDFFFF80021FFFEFFDF000A",
		INIT_37=>X"FFDDFFED00260007FFD800020026FFF3FFDD0015001CFFE3FFEA0021000CFFDB",
		INIT_38=>X"0029FFE5FFDD00220018FFD7FFF1002B0002FFD400080028FFEDFFDD001B001B",
		INIT_39=>X"FFFD0035FFF4FFCE0017002AFFDDFFDE002A0015FFD1FFF60030FFFCFFD1000F",
		INIT_3A=>X"FFC8FFE4003C000AFFC10005003BFFEBFFCB0021002AFFD4FFE100320010FFC9",
		INIT_3B=>X"0047FFD1FFC6003C0028FFBBFFEA00480002FFB8000F0041FFDFFFC8002D002A",
		INIT_3C=>X"FFFD0069FFE7FFA0002F004FFFBDFFC4004F0025FFA9FFF10057FFF7FFAD001D",
		INIT_3D=>X"FF74FFC100930016FF6F000F0085FFCFFF8D004B0059FFA1FFC2006A001FFF92",
		INIT_3E=>X"011BFF47FF3100D80084FF1BFFC000E00002FF30003100B3FFA5FF6F00790068",
		INIT_3F=>X"22A81432FD5FF9B80289033DFD9BFE38023300E0FE08FFBF01B2FFCEFE970082",
		INIT_40=>X"0007FFFCFFFD0007FFF800030002FFF90007FFFBFFFE0006FFF800050000FFFA",
		INIT_41=>X"00050000FFFA0008FFFA00000005FFF80006FFFEFFFB0007FFF900020003FFF8",
		INIT_42=>X"00020003FFF80007FFFCFFFD0007FFF800040001FFF90007FFFBFFFE0006FFF8",
		INIT_43=>X"FFFF0006FFF70005FFFFFFFA0008FFF900000004FFF80006FFFEFFFB0007FFF8",
		INIT_44=>X"FFFC0007FFF800020003FFF80007FFFCFFFD0007FFF800040001FFF90007FFFB",
		INIT_45=>X"FFF90008FFFAFFFF0005FFF70005FFFFFFFA0008FFF900010004FFF80006FFFE",
		INIT_46=>X"FFF80006FFFDFFFC0007FFF800020003FFF80007FFFCFFFD0006FFF800040001",
		INIT_47=>X"FFF800040001FFF90008FFFAFFFF0005FFF70005FFFFFFFA0008FFF900010004",
		INIT_48=>X"FFF900010004FFF80007FFFDFFFC0007FFF800030002FFF80007FFFCFFFD0006",
		INIT_49=>X"FFFBFFFE0006FFF700040000FFF90008FFFAFFFF0005FFF70006FFFFFFFA0008",
		INIT_4A=>X"FFFEFFFB0008FFF900010004FFF80007FFFDFFFC0007FFF800030002FFF80007",
		INIT_4B=>X"0002FFF80008FFFBFFFE0006FFF700050000FFF90008FFFA00000005FFF70006",
		INIT_4C=>X"0005FFF70006FFFEFFFB0008FFF800020004FFF80007FFFDFFFC0007FFF80003",
		INIT_4D=>X"0007FFF700040002FFF80008FFFBFFFE0006FFF700050000FFF90008FFF90000",
		INIT_4E=>X"0008FFF900000005FFF70006FFFEFFFB0008FFF800020003FFF70007FFFCFFFC",
		INIT_4F=>X"0008FFFCFFFD0007FFF700040002FFF80008FFFAFFFE0006FFF700050000FFF9",
		INIT_50=>X"0006FFFFFFF90008FFF900000005FFF70007FFFEFFFB0008FFF800020003FFF7",
		INIT_51=>X"00020003FFF70008FFFCFFFD0007FFF700040001FFF80008FFFAFFFF0006FFF7",
		INIT_52=>X"FFFF0006FFF70006FFFFFFFA0008FFF900010005FFF70007FFFDFFFB0008FFF8",
		INIT_53=>X"FFFB0008FFF700030003FFF70008FFFBFFFD0007FFF700040001FFF80008FFFA",
		INIT_54=>X"FFF80009FFF9FFFF0006FFF60006FFFFFFFA0009FFF800010005FFF70007FFFD",
		INIT_55=>X"FFF60008FFFDFFFB0008FFF700030003FFF70008FFFBFFFD0007FFF600050001",
		INIT_56=>X"FFF600050001FFF80009FFF9FFFF0006FFF60007FFFFFFFA0009FFF800010005",
		INIT_57=>X"FFF800020004FFF60008FFFCFFFB0008FFF700030003FFF70009FFFBFFFD0007",
		INIT_58=>X"FFFAFFFE0007FFF600060000FFF80009FFF900000006FFF60007FFFEFFFA0009",
		INIT_59=>X"FFFEFFFA0009FFF700020004FFF60008FFFCFFFC0009FFF600040002FFF70009",
		INIT_5A=>X"0002FFF70009FFFAFFFE0008FFF500060000FFF8000AFFF800000006FFF60007",
		INIT_5B=>X"0006FFF50008FFFEFFFA000AFFF700020004FFF60009FFFCFFFC0009FFF60004",
		INIT_5C=>X"0009FFF500050002FFF7000AFFF9FFFE0008FFF500060000FFF8000AFFF80000",
		INIT_5D=>X"000AFFF700010006FFF50008FFFDFFFA000AFFF600030004FFF60009FFFBFFFC",
		INIT_5E=>X"000AFFFBFFFC0009FFF500050002FFF6000AFFF9FFFE0008FFF500070000FFF8",
		INIT_5F=>X"0008FFFFFFF8000BFFF700010006FFF40009FFFDFFFA000AFFF600030004FFF5",
		INIT_60=>X"00040004FFF5000AFFFAFFFC0009FFF400060002FFF6000BFFF8FFFF0008FFF4",
		INIT_61=>X"FFFF0008FFF40008FFFFFFF8000BFFF600010006FFF40009FFFCFFFA000BFFF5",
		INIT_62=>X"FFFA000BFFF400040004FFF5000BFFFAFFFC000AFFF400060001FFF6000BFFF8",
		INIT_63=>X"FFF6000CFFF7FFFF0008FFF30009FFFEFFF8000CFFF500020006FFF4000AFFFC",
		INIT_64=>X"FFF3000BFFFBFFFA000CFFF400050004FFF4000CFFF9FFFD000AFFF300070001",
		INIT_65=>X"FFF200080001FFF5000DFFF600000009FFF2000AFFFEFFF8000CFFF500020006",
		INIT_66=>X"FFF400030006FFF2000CFFFBFFFA000CFFF300050004FFF4000DFFF8FFFD000B",
		INIT_67=>X"FFF8FFFD000BFFF100090000FFF5000EFFF500000009FFF2000AFFFEFFF7000D",
		INIT_68=>X"FFFDFFF7000EFFF300040006FFF2000DFFFAFFFA000DFFF200060003FFF3000E",
		INIT_69=>X"0003FFF2000FFFF7FFFD000CFFF0000A0000FFF5000FFFF400010009FFF1000C",
		INIT_6A=>X"0009FFEF000DFFFCFFF7000FFFF200040006FFF1000EFFF9FFFA000EFFF10007",
		INIT_6B=>X"000EFFEF00080003FFF20010FFF5FFFE000CFFEF000B0000FFF40010FFF30001",
		INIT_6C=>X"0011FFF20002000AFFEE000EFFFCFFF70010FFF000050007FFF0000FFFF8FFFA",
		INIT_6D=>X"0011FFF7FFFA0010FFEE00090003FFF10012FFF4FFFE000DFFED000CFFFFFFF3",
		INIT_6E=>X"000EFFFFFFF30013FFF00002000AFFED0010FFFBFFF60012FFEE00060007FFEE",
		INIT_6F=>X"00080007FFED0013FFF6FFFA0011FFEC000B0003FFEF0013FFF3FFFE000EFFEC",
		INIT_70=>X"FFFF000FFFE90010FFFEFFF20015FFEE0003000BFFEB0012FFF9FFF60013FFEC",
		INIT_71=>X"FFF50016FFEA00090007FFEB0016FFF4FFFA0013FFE9000D0002FFEE0016FFF1",
		INIT_72=>X"FFEC0019FFEE00000011FFE70012FFFDFFF10018FFEB0005000CFFE80015FFF8",
		INIT_73=>X"FFE50018FFF6FFF50018FFE6000B0008FFE80019FFF2FFFA0015FFE6000F0002",
		INIT_74=>X"FFE200120002FFEA001DFFEB00000013FFE30016FFFCFFEF001BFFE80006000D",
		INIT_75=>X"FFE30008000FFFE1001DFFF4FFF4001CFFE2000E0008FFE5001DFFEFFFFA0018",
		INIT_76=>X"FFEAFFFA001CFFDC00170001FFE60022FFE600020015FFDE001AFFFAFFED0020",
		INIT_77=>X"FFF8FFEA0027FFDD000B0011FFDB0023FFF0FFF20022FFDB00120009FFE00024",
		INIT_78=>X"000AFFD9002DFFE4FFFA0022FFD3001D0000FFE1002AFFDF00030019FFD60021",
		INIT_79=>X"0020FFCA002CFFF4FFE50031FFD200100014FFD1002DFFEBFFF0002AFFD20018",
		INIT_7A=>X"0038FFC10022000CFFCD003CFFDAFFFA002CFFC50028FFFFFFD90038FFD50006",
		INIT_7B=>X"0051FFC0000B002CFFB40040FFEDFFDC0045FFBF0018001BFFC0003FFFE2FFEC",
		INIT_7C=>X"0067FFCDFFE40057FF9D0037000FFFB4005CFFC4FFFA0040FFA8003DFFFCFFC9",
		INIT_7D=>X"0078FFF4FF9F0093FF8B0019004BFF7D0070FFDCFFC70072FF93002B0029FF9B",
		INIT_7E=>X"00840066FEFD0107FF7EFFC500C7FF21007F001BFF6300C0FF83FFFA007BFF57",
		INIT_7F=>X"30880E06F5D30529FF78FD84035AFD9A0087012FFE0801A0FF7AFF52015BFEBE",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_14,
		DOPADOP=>dopadop_14,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_15: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"C33CCF30CF30CF30CF33CC33CC33CC33CCF30CF30CF30CF30CC33CC33CC33CC3",
		INITP_01=>X"3CC33CC330CF30CF30CF30CC33CC33CC33CC330CF30CF30CF30CF33CC33CC33C",
		INITP_02=>X"C33CC33CC33CCF30CF30CF30CF33CC33CC33CC33CCF30CF30CF30CF33CC33CC3",
		INITP_03=>X"3CC33CC33CC33CC330CF30CF30CF30CC33CC33CC33CC330CF30CF30CF30CC33C",
		INITP_04=>X"F30CC33CC33CC33CC330CF30CF30CF30CF33CC33CC33CC33CCF30CF30CF30CF3",
		INITP_05=>X"0CF30CF33CC33CC33CC33CCF30CF30CF30CF30CC33CC33CC33CC330CF30CF30C",
		INITP_06=>X"F30CF30CF30CC33CC33CC33CC330CF30CF30CF30CC33CC33CC33CC33CCF30CF3",
		INITP_07=>X"0CF30CF30CF30CF33CC33CC33CC33CCF30CF30CF30CF33CC33CC33CC33CC330C",
		INITP_08=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_09=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000",
		INITP_0A=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0B=>X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0C=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_0D=>X"FFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0F=>X"3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_00=>X"0007FFFCFFFD0007FFF800030002FFF90007FFFBFFFE0006FFF800050000FFFA",
		INIT_01=>X"00050000FFFA0008FFFA00000005FFF80006FFFEFFFB0007FFF900020003FFF8",
		INIT_02=>X"00020003FFF80007FFFCFFFD0007FFF800040001FFF90007FFFBFFFE0006FFF8",
		INIT_03=>X"FFFF0006FFF70005FFFFFFFA0008FFF900000004FFF80006FFFEFFFB0007FFF8",
		INIT_04=>X"FFFC0007FFF800020003FFF80007FFFCFFFD0007FFF800040001FFF90007FFFB",
		INIT_05=>X"FFF90008FFFAFFFF0005FFF70005FFFFFFFA0008FFF900010004FFF80006FFFE",
		INIT_06=>X"FFF80006FFFDFFFC0007FFF800020003FFF80007FFFCFFFD0006FFF800040001",
		INIT_07=>X"FFF800040001FFF90008FFFAFFFF0005FFF70005FFFFFFFA0008FFF900010004",
		INIT_08=>X"FFF900010004FFF80007FFFDFFFC0007FFF800030002FFF80007FFFCFFFD0006",
		INIT_09=>X"FFFBFFFE0006FFF700040000FFF90008FFFAFFFF0005FFF70006FFFFFFFA0008",
		INIT_0A=>X"FFFEFFFB0008FFF900010004FFF80007FFFDFFFC0007FFF800030002FFF80007",
		INIT_0B=>X"0002FFF80008FFFBFFFE0006FFF700050000FFF90008FFFA00000005FFF70006",
		INIT_0C=>X"0005FFF70006FFFEFFFB0008FFF800020004FFF80007FFFDFFFC0007FFF80003",
		INIT_0D=>X"0007FFF700040002FFF80008FFFBFFFE0006FFF700050000FFF90008FFF90000",
		INIT_0E=>X"0008FFF900000005FFF70006FFFEFFFB0008FFF800020003FFF70007FFFCFFFC",
		INIT_0F=>X"0008FFFCFFFD0007FFF700040002FFF80008FFFAFFFE0006FFF700050000FFF9",
		INIT_10=>X"0006FFFFFFF90008FFF900000005FFF70007FFFEFFFB0008FFF800020003FFF7",
		INIT_11=>X"00020003FFF70008FFFCFFFD0007FFF700040001FFF80008FFFAFFFF0006FFF7",
		INIT_12=>X"FFFF0006FFF70006FFFFFFFA0008FFF900010005FFF70007FFFDFFFB0008FFF8",
		INIT_13=>X"FFFB0008FFF700030003FFF70008FFFBFFFD0007FFF700040001FFF80008FFFA",
		INIT_14=>X"FFF80009FFF9FFFF0006FFF60006FFFFFFFA0009FFF800010005FFF70007FFFD",
		INIT_15=>X"FFF60008FFFDFFFB0008FFF700030003FFF70008FFFBFFFD0007FFF600050001",
		INIT_16=>X"FFF600050001FFF80009FFF9FFFF0006FFF60007FFFFFFFA0009FFF800010005",
		INIT_17=>X"FFF800020004FFF60008FFFCFFFB0008FFF700030003FFF70009FFFBFFFD0007",
		INIT_18=>X"FFFAFFFE0007FFF600060000FFF80009FFF900000006FFF60007FFFEFFFA0009",
		INIT_19=>X"FFFEFFFA0009FFF700020004FFF60008FFFCFFFC0009FFF600040002FFF70009",
		INIT_1A=>X"0002FFF70009FFFAFFFE0008FFF500060000FFF8000AFFF800000006FFF60007",
		INIT_1B=>X"0006FFF50008FFFEFFFA000AFFF700020004FFF60009FFFCFFFC0009FFF60004",
		INIT_1C=>X"0009FFF500050002FFF7000AFFF9FFFE0008FFF500060000FFF8000AFFF80000",
		INIT_1D=>X"000AFFF700010006FFF50008FFFDFFFA000AFFF600030004FFF60009FFFBFFFC",
		INIT_1E=>X"000AFFFBFFFC0009FFF500050002FFF6000AFFF9FFFE0008FFF500070000FFF8",
		INIT_1F=>X"0008FFFFFFF8000BFFF700010006FFF40009FFFDFFFA000AFFF600030004FFF5",
		INIT_20=>X"00040004FFF5000AFFFAFFFC0009FFF400060002FFF6000BFFF8FFFF0008FFF4",
		INIT_21=>X"FFFF0008FFF40008FFFFFFF8000BFFF600010006FFF40009FFFCFFFA000BFFF5",
		INIT_22=>X"FFFA000BFFF400040004FFF5000BFFFAFFFC000AFFF400060001FFF6000BFFF8",
		INIT_23=>X"FFF6000CFFF7FFFF0008FFF30009FFFEFFF8000CFFF500020006FFF4000AFFFC",
		INIT_24=>X"FFF3000BFFFBFFFA000CFFF400050004FFF4000CFFF9FFFD000AFFF300070001",
		INIT_25=>X"FFF200080001FFF5000DFFF600000009FFF2000AFFFEFFF8000CFFF500020006",
		INIT_26=>X"FFF400030006FFF2000CFFFBFFFA000CFFF300050004FFF4000DFFF8FFFD000B",
		INIT_27=>X"FFF8FFFD000BFFF100090000FFF5000EFFF500000009FFF2000AFFFEFFF7000D",
		INIT_28=>X"FFFDFFF7000EFFF300040006FFF2000DFFFAFFFA000DFFF200060003FFF3000E",
		INIT_29=>X"0003FFF2000FFFF7FFFD000CFFF0000A0000FFF5000FFFF400010009FFF1000C",
		INIT_2A=>X"0009FFEF000DFFFCFFF7000FFFF200040006FFF1000EFFF9FFFA000EFFF10007",
		INIT_2B=>X"000EFFEF00080003FFF20010FFF5FFFE000CFFEF000B0000FFF40010FFF30001",
		INIT_2C=>X"0011FFF20002000AFFEE000EFFFCFFF70010FFF000050007FFF0000FFFF8FFFA",
		INIT_2D=>X"0011FFF7FFFA0010FFEE00090003FFF10012FFF4FFFE000DFFED000CFFFFFFF3",
		INIT_2E=>X"000EFFFFFFF30013FFF00002000AFFED0010FFFBFFF60012FFEE00060007FFEE",
		INIT_2F=>X"00080007FFED0013FFF6FFFA0011FFEC000B0003FFEF0013FFF3FFFE000EFFEC",
		INIT_30=>X"FFFF000FFFE90010FFFEFFF20015FFEE0003000BFFEB0012FFF9FFF60013FFEC",
		INIT_31=>X"FFF50016FFEA00090007FFEB0016FFF4FFFA0013FFE9000D0002FFEE0016FFF1",
		INIT_32=>X"FFEC0019FFEE00000011FFE70012FFFDFFF10018FFEB0005000CFFE80015FFF8",
		INIT_33=>X"FFE50018FFF6FFF50018FFE6000B0008FFE80019FFF2FFFA0015FFE6000F0002",
		INIT_34=>X"FFE200120002FFEA001DFFEB00000013FFE30016FFFCFFEF001BFFE80006000D",
		INIT_35=>X"FFE30008000FFFE1001DFFF4FFF4001CFFE2000E0008FFE5001DFFEFFFFA0018",
		INIT_36=>X"FFEAFFFA001CFFDC00170001FFE60022FFE600020015FFDE001AFFFAFFED0020",
		INIT_37=>X"FFF8FFEA0027FFDD000B0011FFDB0023FFF0FFF20022FFDB00120009FFE00024",
		INIT_38=>X"000AFFD9002DFFE4FFFA0022FFD3001D0000FFE1002AFFDF00030019FFD60021",
		INIT_39=>X"0020FFCA002CFFF4FFE50031FFD200100014FFD1002DFFEBFFF0002AFFD20018",
		INIT_3A=>X"0038FFC10022000CFFCD003CFFDAFFFA002CFFC50028FFFFFFD90038FFD50006",
		INIT_3B=>X"0051FFC0000B002CFFB40040FFEDFFDC0045FFBF0018001BFFC0003FFFE2FFEC",
		INIT_3C=>X"0067FFCDFFE40057FF9D0037000FFFB4005CFFC4FFFA0040FFA8003DFFFCFFC9",
		INIT_3D=>X"0078FFF4FF9F0093FF8B0019004BFF7D0070FFDCFFC70072FF93002B0029FF9B",
		INIT_3E=>X"00840066FEFD0107FF7EFFC500C7FF21007F001BFF6300C0FF83FFFA007BFF57",
		INIT_3F=>X"30880E06F5D30529FF78FD84035AFD9A0087012FFE0801A0FF7AFF52015BFEBE",
		INIT_40=>X"0007000700070007000700070007000700070007000700070007000700070007",
		INIT_41=>X"0007000700070007000700070007000700070007000700070007000700070007",
		INIT_42=>X"0006000700070007000700070007000700070007000700070007000700070007",
		INIT_43=>X"0006000600060006000600060006000600060006000600060006000600060006",
		INIT_44=>X"0005000500050005000500050005000500050005000500050005000600060006",
		INIT_45=>X"0004000400040004000400040004000400040004000400040005000500050005",
		INIT_46=>X"0002000300030003000300030003000300030003000300030003000300040004",
		INIT_47=>X"0001000100010001000100020002000200020002000200020002000200020002",
		INIT_48=>X"0000000000000000000000000000000000000000000100010001000100010001",
		INIT_49=>X"FFFEFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000",
		INIT_4A=>X"FFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFE",
		INIT_4B=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFD",
		INIT_4C=>X"FFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFB",
		INIT_4D=>X"FFF9FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFA",
		INIT_4E=>X"FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_4F=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_50=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_51=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_52=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_53=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_54=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_55=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7",
		INIT_56=>X"FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_57=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_58=>X"FFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFA",
		INIT_59=>X"FFFDFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFC",
		INIT_5A=>X"FFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFD",
		INIT_5B=>X"0001000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_5C=>X"0002000200020002000200020002000200010001000100010001000100010001",
		INIT_5D=>X"0004000400040004000400040003000300030003000300030003000300030002",
		INIT_5E=>X"0006000600060006000500050005000500050005000500050005000400040004",
		INIT_5F=>X"0008000700070007000700070007000700070007000600060006000600060006",
		INIT_60=>X"0009000900090009000900090008000800080008000800080008000800080008",
		INIT_61=>X"000A000A000A000A000A000A000A000A000A000A000900090009000900090009",
		INIT_62=>X"000B000B000B000B000B000B000B000B000B000B000B000B000B000A000A000A",
		INIT_63=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000B000B000B",
		INIT_64=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C",
		INIT_65=>X"000D000D000D000D000D000D000D000D000D000D000D000D000D000D000C000C",
		INIT_66=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000C000D000D",
		INIT_67=>X"000B000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C",
		INIT_68=>X"000A000A000A000B000B000B000B000B000B000B000B000B000B000B000B000B",
		INIT_69=>X"0009000900090009000900090009000A000A000A000A000A000A000A000A000A",
		INIT_6A=>X"0007000700070007000700070008000800080008000800080008000800090009",
		INIT_6B=>X"0004000500050005000500050005000600060006000600060006000600070007",
		INIT_6C=>X"0002000200020002000200030003000300030003000300040004000400040004",
		INIT_6D=>X"FFFFFFFFFFFFFFFFFFFF00000000000000000000000100010001000100010001",
		INIT_6E=>X"FFFBFFFBFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFE",
		INIT_6F=>X"FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFB",
		INIT_70=>X"FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7",
		INIT_71=>X"FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3",
		INIT_72=>X"FFEBFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEFFFEFFFEFFFEF",
		INIT_73=>X"FFE7FFE7FFE8FFE8FFE8FFE9FFE9FFE9FFE9FFEAFFEAFFEAFFEAFFEBFFEBFFEB",
		INIT_74=>X"FFE3FFE3FFE4FFE4FFE4FFE4FFE5FFE5FFE5FFE5FFE6FFE6FFE6FFE6FFE7FFE7",
		INIT_75=>X"FFDFFFDFFFDFFFE0FFE0FFE0FFE0FFE1FFE1FFE1FFE1FFE2FFE2FFE2FFE3FFE3",
		INIT_76=>X"FFDBFFDBFFDBFFDCFFDCFFDCFFDCFFDDFFDDFFDDFFDDFFDEFFDEFFDEFFDEFFDF",
		INIT_77=>X"FFD7FFD8FFD8FFD8FFD8FFD8FFD9FFD9FFD9FFD9FFDAFFDAFFDAFFDAFFDBFFDB",
		INIT_78=>X"FFD4FFD4FFD4FFD4FFD5FFD5FFD5FFD5FFD6FFD6FFD6FFD6FFD6FFD7FFD7FFD7",
		INIT_79=>X"FFD1FFD1FFD1FFD1FFD1FFD2FFD2FFD2FFD2FFD2FFD3FFD3FFD3FFD3FFD3FFD4",
		INIT_7A=>X"FFCEFFCEFFCEFFCEFFCFFFCFFFCFFFCFFFCFFFCFFFD0FFD0FFD0FFD0FFD0FFD1",
		INIT_7B=>X"FFCCFFCCFFCCFFCCFFCCFFCCFFCDFFCDFFCDFFCDFFCDFFCDFFCDFFCEFFCEFFCE",
		INIT_7C=>X"FFCAFFCAFFCAFFCAFFCAFFCAFFCBFFCBFFCBFFCBFFCBFFCBFFCBFFCBFFCBFFCC",
		INIT_7D=>X"FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFCAFFCAFFCAFFCA",
		INIT_7E=>X"FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC9",
		INIT_7F=>X"3FC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_15,
		DOPADOP=>dopadop_15,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
end arch;
