library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity filter_table is
	port(
		clk:  in  std_logic;
		addr: in  std_logic_vector(14 downto 0);
		data: out signed(17 downto 0)
	);
end filter_table;

architecture arch of filter_table is
	signal addr_d:  std_logic_vector(14 downto 11);
	signal addrardaddr:   std_logic_vector(15 downto 0);
	signal doado_00:  std_logic_vector(31 downto 0);
	signal dopadop_00: std_logic_vector(3 downto 0);
	signal doado_01:  std_logic_vector(31 downto 0);
	signal dopadop_01: std_logic_vector(3 downto 0);
	signal doado_02:  std_logic_vector(31 downto 0);
	signal dopadop_02: std_logic_vector(3 downto 0);
	signal doado_03:  std_logic_vector(31 downto 0);
	signal dopadop_03: std_logic_vector(3 downto 0);
	signal doado_04:  std_logic_vector(31 downto 0);
	signal dopadop_04: std_logic_vector(3 downto 0);
	signal doado_05:  std_logic_vector(31 downto 0);
	signal dopadop_05: std_logic_vector(3 downto 0);
	signal doado_06:  std_logic_vector(31 downto 0);
	signal dopadop_06: std_logic_vector(3 downto 0);
	signal doado_07:  std_logic_vector(31 downto 0);
	signal dopadop_07: std_logic_vector(3 downto 0);
	signal doado_08:  std_logic_vector(31 downto 0);
	signal dopadop_08: std_logic_vector(3 downto 0);
	signal doado_09:  std_logic_vector(31 downto 0);
	signal dopadop_09: std_logic_vector(3 downto 0);
	signal doado_10:  std_logic_vector(31 downto 0);
	signal dopadop_10: std_logic_vector(3 downto 0);
	signal doado_11:  std_logic_vector(31 downto 0);
	signal dopadop_11: std_logic_vector(3 downto 0);
	signal doado_12:  std_logic_vector(31 downto 0);
	signal dopadop_12: std_logic_vector(3 downto 0);
	signal doado_13:  std_logic_vector(31 downto 0);
	signal dopadop_13: std_logic_vector(3 downto 0);
	signal doado_14:  std_logic_vector(31 downto 0);
	signal dopadop_14: std_logic_vector(3 downto 0);
	signal doado_15:  std_logic_vector(31 downto 0);
	signal dopadop_15: std_logic_vector(3 downto 0);
begin
	addrardaddr(15)<='1';
	addrardaddr(14 downto 4)<=addr(10 downto 0);
	addrardaddr(3 downto 0)<=b"0000";
	process(clk)
	begin
		if (rising_edge(clk)) then
			addr_d<=addr(14 downto 11);
		end if;
	end process;
	with addr_d select data(15 downto 0)<=
		signed(doado_00(15 downto 0)) when b"0000",
		signed(doado_01(15 downto 0)) when b"0001",
		signed(doado_02(15 downto 0)) when b"0010",
		signed(doado_03(15 downto 0)) when b"0011",
		signed(doado_04(15 downto 0)) when b"0100",
		signed(doado_05(15 downto 0)) when b"0101",
		signed(doado_06(15 downto 0)) when b"0110",
		signed(doado_07(15 downto 0)) when b"0111",
		signed(doado_08(15 downto 0)) when b"1000",
		signed(doado_09(15 downto 0)) when b"1001",
		signed(doado_10(15 downto 0)) when b"1010",
		signed(doado_11(15 downto 0)) when b"1011",
		signed(doado_12(15 downto 0)) when b"1100",
		signed(doado_13(15 downto 0)) when b"1101",
		signed(doado_14(15 downto 0)) when b"1110",
		signed(doado_15(15 downto 0)) when others;
	with addr_d select data(17 downto 16)<=
		signed(dopadop_00(1 downto 0)) when b"0000",
		signed(dopadop_01(1 downto 0)) when b"0001",
		signed(dopadop_02(1 downto 0)) when b"0010",
		signed(dopadop_03(1 downto 0)) when b"0011",
		signed(dopadop_04(1 downto 0)) when b"0100",
		signed(dopadop_05(1 downto 0)) when b"0101",
		signed(dopadop_06(1 downto 0)) when b"0110",
		signed(dopadop_07(1 downto 0)) when b"0111",
		signed(dopadop_08(1 downto 0)) when b"1000",
		signed(dopadop_09(1 downto 0)) when b"1001",
		signed(dopadop_10(1 downto 0)) when b"1010",
		signed(dopadop_11(1 downto 0)) when b"1011",
		signed(dopadop_12(1 downto 0)) when b"1100",
		signed(dopadop_13(1 downto 0)) when b"1101",
		signed(dopadop_14(1 downto 0)) when b"1110",
		signed(dopadop_15(1 downto 0)) when others;
	mem_00: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02=>X"FFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000",
		INITP_03=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_04=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_05=>X"0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF",
		INITP_06=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_08=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_09=>X"FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000",
		INITP_0A=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0B=>X"000000000000000000000000000000000000000000000000000FFFFFFFFFFFFF",
		INITP_0C=>X"FFFFFFFFFFFFC000000000000000000000000000000000000000000000000000",
		INITP_0D=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0E=>X"00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0F=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_00=>X"002F002F002F002F002F002F002F002F002F002F002F002F002F002F002F0030",
		INIT_01=>X"002F002F002F002F002F002F002F002F002F002F002F002F002F002F002F002F",
		INIT_02=>X"002E002E002E002E002E002E002E002F002F002F002F002F002F002F002F002F",
		INIT_03=>X"002D002D002D002D002D002D002E002E002E002E002E002E002E002E002E002E",
		INIT_04=>X"002C002C002C002C002C002C002C002C002D002D002D002D002D002D002D002D",
		INIT_05=>X"002A002A002A002B002B002B002B002B002B002B002B002B002B002C002C002C",
		INIT_06=>X"0028002800290029002900290029002900290029002A002A002A002A002A002A",
		INIT_07=>X"0026002600270027002700270027002700270027002800280028002800280028",
		INIT_08=>X"0024002400240024002500250025002500250025002500260026002600260026",
		INIT_09=>X"0021002200220022002200220022002300230023002300230023002300240024",
		INIT_0A=>X"001F001F001F001F001F00200020002000200020002000210021002100210021",
		INIT_0B=>X"001C001C001C001C001D001D001D001D001D001E001E001E001E001E001E001F",
		INIT_0C=>X"001900190019001A001A001A001A001A001A001B001B001B001B001B001C001C",
		INIT_0D=>X"0016001600160017001700170017001700170018001800180018001800190019",
		INIT_0E=>X"0013001300130013001400140014001400140015001500150015001500160016",
		INIT_0F=>X"0010001000100010001000110011001100110011001200120012001200120013",
		INIT_10=>X"000D000D000D000D000D000E000E000E000E000E000F000F000F000F000F0010",
		INIT_11=>X"0009000A000A000A000A000A000B000B000B000B000B000C000C000C000C000C",
		INIT_12=>X"0006000700070007000700070008000800080008000800080009000900090009",
		INIT_13=>X"0003000400040004000400040005000500050005000500050006000600060006",
		INIT_14=>X"0001000100010001000100010002000200020002000200030003000300030003",
		INIT_15=>X"FFFEFFFEFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000",
		INIT_16=>X"FFFBFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFE",
		INIT_17=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFB",
		INIT_18=>X"FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9",
		INIT_19=>X"FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_1A=>X"FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5",
		INIT_1B=>X"FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3",
		INIT_1C=>X"FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2FFF2FFF2FFF2",
		INIT_1D=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1",
		INIT_1E=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_1F=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_20=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_21=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_22=>X"FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_23=>X"FFF2FFF2FFF2FFF2FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1",
		INIT_24=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2",
		INIT_25=>X"FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF3FFF3FFF3",
		INIT_26=>X"FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5",
		INIT_27=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_28=>X"FFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9",
		INIT_29=>X"FFFEFFFDFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFB",
		INIT_2A=>X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFE",
		INIT_2B=>X"0003000300030003000200020002000200020001000100010001000100010000",
		INIT_2C=>X"0006000600060005000500050005000500050004000400040004000400030003",
		INIT_2D=>X"0009000900090008000800080008000800080007000700070007000700060006",
		INIT_2E=>X"000C000C000C000C000B000B000B000B000B000A000A000A000A000A00090009",
		INIT_2F=>X"000F000F000F000F000F000E000E000E000E000E000D000D000D000D000D000C",
		INIT_30=>X"0012001200120012001200110011001100110011001000100010001000100010",
		INIT_31=>X"0016001500150015001500150014001400140014001400130013001300130013",
		INIT_32=>X"0019001800180018001800180017001700170017001700170016001600160016",
		INIT_33=>X"001C001B001B001B001B001B001A001A001A001A001A001A0019001900190019",
		INIT_34=>X"001E001E001E001E001E001E001D001D001D001D001D001C001C001C001C001C",
		INIT_35=>X"0021002100210021002000200020002000200020001F001F001F001F001F001F",
		INIT_36=>X"0024002300230023002300230023002300220022002200220022002200210021",
		INIT_37=>X"0026002600260026002500250025002500250025002500240024002400240024",
		INIT_38=>X"0028002800280028002800270027002700270027002700270027002600260026",
		INIT_39=>X"002A002A002A002A002A00290029002900290029002900290029002800280028",
		INIT_3A=>X"002C002C002B002B002B002B002B002B002B002B002B002B002A002A002A002A",
		INIT_3B=>X"002D002D002D002D002D002D002D002C002C002C002C002C002C002C002C002C",
		INIT_3C=>X"002E002E002E002E002E002E002E002E002E002D002D002D002D002D002D002D",
		INIT_3D=>X"002F002F002F002F002F002F002F002F002E002E002E002E002E002E002E002E",
		INIT_3E=>X"002F002F002F002F002F002F002F002F002F002F002F002F002F002F002F002F",
		INIT_3F=>X"002F002F002F002F002F002F002F002F002F002F002F002F002F002F002F002F",
		INIT_40=>X"004F004F004F004F004F004F004F004F004F004F004F004F004F004F004F0050",
		INIT_41=>X"004D004D004D004D004D004D004E004E004E004E004E004E004E004F004F004F",
		INIT_42=>X"00490049004A004A004A004A004B004B004B004B004B004C004C004C004C004C",
		INIT_43=>X"0044004400450045004500460046004600470047004700480048004800480049",
		INIT_44=>X"003E003E003F003F004000400040004100410041004200420043004300430044",
		INIT_45=>X"003700370038003800390039003A003A003A003B003B003C003C003D003D003D",
		INIT_46=>X"002F002F00300031003100320032003200330033003400340035003500360036",
		INIT_47=>X"002700270028002800290029002A002A002B002B002C002C002D002D002E002E",
		INIT_48=>X"001E001F001F0020002000210021002200220023002300240025002500260026",
		INIT_49=>X"00160016001700170018001800190019001A001A001B001B001C001C001D001E",
		INIT_4A=>X"000D000E000E000F000F00100010001100110012001200130013001400150015",
		INIT_4B=>X"000600060007000700070008000800090009000A000A000B000B000C000C000D",
		INIT_4C=>X"FFFFFFFFFFFF0000000000010001000200020002000300030004000400050005",
		INIT_4D=>X"FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFDFFFDFFFDFFFEFFFE",
		INIT_4E=>X"FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF8FFF8",
		INIT_4F=>X"FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2FFF3FFF3FFF3",
		INIT_50=>X"FFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEFFFEFFFF0",
		INIT_51=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFED",
		INIT_52=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_53=>X"FFEDFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_54=>X"FFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFED",
		INIT_55=>X"FFF1FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEF",
		INIT_56=>X"FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF1",
		INIT_57=>X"FFF9FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5",
		INIT_58=>X"FFFDFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFF9FFF9FFF9",
		INIT_59=>X"000100010000000000000000FFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFDFFFD",
		INIT_5A=>X"0005000500040004000400040003000300030003000200020002000200010001",
		INIT_5B=>X"0008000800080008000800070007000700070006000600060006000600050005",
		INIT_5C=>X"000B000B000B000B000B000A000A000A000A000A000A00090009000900090009",
		INIT_5D=>X"000E000D000D000D000D000D000D000D000D000C000C000C000C000C000C000B",
		INIT_5E=>X"000F000F000F000F000F000F000F000E000E000E000E000E000E000E000E000E",
		INIT_5F=>X"000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F",
		INIT_60=>X"000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F0010",
		INIT_61=>X"000E000E000E000E000E000E000E000E000F000F000F000F000F000F000F000F",
		INIT_62=>X"000C000C000C000C000C000C000D000D000D000D000D000D000D000D000E000E",
		INIT_63=>X"0009000900090009000A000A000A000A000A000A000B000B000B000B000B000B",
		INIT_64=>X"0005000600060006000600060007000700070007000800080008000800080009",
		INIT_65=>X"0001000200020002000200030003000300030004000400040004000500050005",
		INIT_66=>X"FFFDFFFEFFFEFFFEFFFEFFFFFFFFFFFFFFFF0000000000000000000100010001",
		INIT_67=>X"FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFD",
		INIT_68=>X"FFF5FFF5FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9",
		INIT_69=>X"FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5",
		INIT_6A=>X"FFEFFFEFFFEFFFEFFFEFFFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF1",
		INIT_6B=>X"FFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEF",
		INIT_6C=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEDFFED",
		INIT_6D=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_6E=>X"FFEDFFEDFFEDFFEDFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_6F=>X"FFEFFFEFFFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFED",
		INIT_70=>X"FFF3FFF3FFF2FFF2FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFF0",
		INIT_71=>X"FFF8FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF3",
		INIT_72=>X"FFFEFFFDFFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8",
		INIT_73=>X"000500040004000300030002000200020001000100000000FFFFFFFFFFFFFFFE",
		INIT_74=>X"000C000C000B000B000A000A0009000900080008000700070007000600060005",
		INIT_75=>X"0015001400130013001200120011001100100010000F000F000E000E000D000D",
		INIT_76=>X"001D001C001C001B001B001A001A001900190018001800170017001600160015",
		INIT_77=>X"002600250025002400230023002200220021002100200020001F001F001E001E",
		INIT_78=>X"002E002D002D002C002C002B002B002A002A0029002900280028002700270026",
		INIT_79=>X"0036003500350034003400330033003200320032003100310030002F002F002E",
		INIT_7A=>X"003D003D003C003C003B003B003A003A003A0039003900380038003700370036",
		INIT_7B=>X"00430043004300420042004100410041004000400040003F003F003E003E003D",
		INIT_7C=>X"0048004800480048004700470047004600460046004500450045004400440044",
		INIT_7D=>X"004C004C004C004C004B004B004B004B004B004A004A004A004A004900490049",
		INIT_7E=>X"004F004F004E004E004E004E004E004E004E004D004D004D004D004D004D004C",
		INIT_7F=>X"004F004F004F004F004F004F004F004F004F004F004F004F004F004F004F004F",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_00,
		DOPADOP=>dopadop_00,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_01: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01=>X"FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000",
		INITP_02=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_03=>X"000000000000000000000000000000000000000000000000000FFFFFFFFFFFFF",
		INITP_04=>X"FFFFFFFFFFFFC000000000000000000000000000000000000000000000000000",
		INITP_05=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_06=>X"00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_08=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_09=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000",
		INITP_0A=>X"0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFF",
		INITP_0B=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000",
		INITP_0C=>X"000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0D=>X"FFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000",
		INITP_0E=>X"000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0F=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_00=>X"004F004F004F004F004F004F004F004F004F004F004F004F004F004F004F0050",
		INIT_01=>X"004D004D004D004D004D004D004E004E004E004E004E004E004E004F004F004F",
		INIT_02=>X"00490049004A004A004A004A004B004B004B004B004B004C004C004C004C004C",
		INIT_03=>X"0044004400450045004500460046004600470047004700480048004800480049",
		INIT_04=>X"003E003E003F003F004000400040004100410041004200420043004300430044",
		INIT_05=>X"003700370038003800390039003A003A003A003B003B003C003C003D003D003D",
		INIT_06=>X"002F002F00300031003100320032003200330033003400340035003500360036",
		INIT_07=>X"002700270028002800290029002A002A002B002B002C002C002D002D002E002E",
		INIT_08=>X"001E001F001F0020002000210021002200220023002300240025002500260026",
		INIT_09=>X"00160016001700170018001800190019001A001A001B001B001C001C001D001E",
		INIT_0A=>X"000D000E000E000F000F00100010001100110012001200130013001400150015",
		INIT_0B=>X"000600060007000700070008000800090009000A000A000B000B000C000C000D",
		INIT_0C=>X"FFFFFFFFFFFF0000000000010001000200020002000300030004000400050005",
		INIT_0D=>X"FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFDFFFDFFFDFFFEFFFE",
		INIT_0E=>X"FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF8FFF8",
		INIT_0F=>X"FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2FFF3FFF3FFF3",
		INIT_10=>X"FFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEFFFEFFFF0",
		INIT_11=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFED",
		INIT_12=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_13=>X"FFEDFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_14=>X"FFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFED",
		INIT_15=>X"FFF1FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEF",
		INIT_16=>X"FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF1",
		INIT_17=>X"FFF9FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5",
		INIT_18=>X"FFFDFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFF9FFF9FFF9",
		INIT_19=>X"000100010000000000000000FFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFDFFFD",
		INIT_1A=>X"0005000500040004000400040003000300030003000200020002000200010001",
		INIT_1B=>X"0008000800080008000800070007000700070006000600060006000600050005",
		INIT_1C=>X"000B000B000B000B000B000A000A000A000A000A000A00090009000900090009",
		INIT_1D=>X"000E000D000D000D000D000D000D000D000D000C000C000C000C000C000C000B",
		INIT_1E=>X"000F000F000F000F000F000F000F000E000E000E000E000E000E000E000E000E",
		INIT_1F=>X"000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F",
		INIT_20=>X"000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F0010",
		INIT_21=>X"000E000E000E000E000E000E000E000E000F000F000F000F000F000F000F000F",
		INIT_22=>X"000C000C000C000C000C000C000D000D000D000D000D000D000D000D000E000E",
		INIT_23=>X"0009000900090009000A000A000A000A000A000A000B000B000B000B000B000B",
		INIT_24=>X"0005000600060006000600060007000700070007000800080008000800080009",
		INIT_25=>X"0001000200020002000200030003000300030004000400040004000500050005",
		INIT_26=>X"FFFDFFFEFFFEFFFEFFFEFFFFFFFFFFFFFFFF0000000000000000000100010001",
		INIT_27=>X"FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFD",
		INIT_28=>X"FFF5FFF5FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9",
		INIT_29=>X"FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5",
		INIT_2A=>X"FFEFFFEFFFEFFFEFFFEFFFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF1",
		INIT_2B=>X"FFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEF",
		INIT_2C=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEDFFED",
		INIT_2D=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_2E=>X"FFEDFFEDFFEDFFEDFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_2F=>X"FFEFFFEFFFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFED",
		INIT_30=>X"FFF3FFF3FFF2FFF2FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFF0",
		INIT_31=>X"FFF8FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF3",
		INIT_32=>X"FFFEFFFDFFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8",
		INIT_33=>X"000500040004000300030002000200020001000100000000FFFFFFFFFFFFFFFE",
		INIT_34=>X"000C000C000B000B000A000A0009000900080008000700070007000600060005",
		INIT_35=>X"0015001400130013001200120011001100100010000F000F000E000E000D000D",
		INIT_36=>X"001D001C001C001B001B001A001A001900190018001800170017001600160015",
		INIT_37=>X"002600250025002400230023002200220021002100200020001F001F001E001E",
		INIT_38=>X"002E002D002D002C002C002B002B002A002A0029002900280028002700270026",
		INIT_39=>X"0036003500350034003400330033003200320032003100310030002F002F002E",
		INIT_3A=>X"003D003D003C003C003B003B003A003A003A0039003900380038003700370036",
		INIT_3B=>X"00430043004300420042004100410041004000400040003F003F003E003E003D",
		INIT_3C=>X"0048004800480048004700470047004600460046004500450045004400440044",
		INIT_3D=>X"004C004C004C004C004B004B004B004B004B004A004A004A004A004900490049",
		INIT_3E=>X"004F004F004E004E004E004E004E004E004E004D004D004D004D004D004D004C",
		INIT_3F=>X"004F004F004F004F004F004F004F004F004F004F004F004F004F004F004F004F",
		INIT_40=>X"006E006E006E006E006E006F006F006F006F006F006F006F006F006F006F0070",
		INIT_41=>X"00680068006900690069006A006A006B006B006B006C006C006C006D006D006D",
		INIT_42=>X"005E005E005F0060006100610062006200630064006400650065006600670067",
		INIT_43=>X"00510052005300530054005500560057005800580059005A005B005C005C005D",
		INIT_44=>X"004200430044004500460047004800490049004A004B004C004D004E004F0050",
		INIT_45=>X"003100320033003400350036003700380039003B003C003D003E003F00400041",
		INIT_46=>X"002000210022002400250026002700280029002A002B002C002D002E002F0030",
		INIT_47=>X"0010001100120013001400150016001700180019001A001B001C001D001E001F",
		INIT_48=>X"000200030004000500060006000700080009000A000B000C000D000E000F000F",
		INIT_49=>X"FFF6FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFCFFFDFFFDFFFEFFFF000000010001",
		INIT_4A=>X"FFEDFFEEFFEEFFEFFFEFFFF0FFF0FFF1FFF1FFF2FFF3FFF3FFF4FFF4FFF5FFF6",
		INIT_4B=>X"FFE8FFE8FFE8FFE9FFE9FFE9FFEAFFEAFFEAFFEBFFEBFFEBFFECFFECFFEDFFED",
		INIT_4C=>X"FFE5FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE7FFE7FFE7FFE7FFE7FFE8",
		INIT_4D=>X"FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE5FFE5FFE5FFE5FFE5FFE5FFE5",
		INIT_4E=>X"FFEAFFE9FFE9FFE9FFE9FFE8FFE8FFE8FFE8FFE7FFE7FFE7FFE7FFE7FFE7FFE6",
		INIT_4F=>X"FFEFFFEFFFEEFFEEFFEEFFEDFFEDFFEDFFECFFECFFECFFEBFFEBFFEBFFEAFFEA",
		INIT_50=>X"FFF6FFF5FFF5FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF2FFF1FFF1FFF0FFF0FFF0",
		INIT_51=>X"FFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF7FFF7FFF6",
		INIT_52=>X"00040004000300030002000200010001000100000000FFFFFFFFFFFEFFFEFFFD",
		INIT_53=>X"000A000A00090009000900080008000700070007000600060006000500050004",
		INIT_54=>X"000E000E000E000E000D000D000D000D000C000C000C000B000B000B000B000A",
		INIT_55=>X"0011001100110010001000100010001000100010000F000F000F000F000F000E",
		INIT_56=>X"0011001100110011001100110011001100110011001100110011001100110011",
		INIT_57=>X"0010001000100010001000100010001100110011001100110011001100110011",
		INIT_58=>X"000C000D000D000D000D000E000E000E000E000E000F000F000F000F000F0010",
		INIT_59=>X"000800080008000900090009000A000A000A000A000B000B000B000C000C000C",
		INIT_5A=>X"0002000300030003000400040004000500050005000600060006000700070007",
		INIT_5B=>X"FFFDFFFDFFFDFFFEFFFEFFFEFFFFFFFFFFFF0000000000010001000100020002",
		INIT_5C=>X"FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFC",
		INIT_5D=>X"FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_5E=>X"FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3FFF3",
		INIT_5F=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_60=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_61=>X"FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF0",
		INIT_62=>X"FFF7FFF7FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3",
		INIT_63=>X"FFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF7FFF7",
		INIT_64=>X"000200010001000100000000FFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFC",
		INIT_65=>X"0007000700060006000600050005000500040004000400030003000300020002",
		INIT_66=>X"000C000C000B000B000B000A000A000A000A0009000900090008000800080007",
		INIT_67=>X"000F000F000F000F000F000E000E000E000E000E000D000D000D000D000C000C",
		INIT_68=>X"0011001100110011001100110011001100100010001000100010001000100010",
		INIT_69=>X"0011001100110011001100110011001100110011001100110011001100110011",
		INIT_6A=>X"000F000F000F000F000F00100010001000100010001000100011001100110011",
		INIT_6B=>X"000B000B000B000B000C000C000C000D000D000D000D000E000E000E000E000E",
		INIT_6C=>X"0005000500060006000600070007000700080008000900090009000A000A000A",
		INIT_6D=>X"FFFEFFFEFFFFFFFF000000000001000100010002000200030003000400040004",
		INIT_6E=>X"FFF7FFF7FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFD",
		INIT_6F=>X"FFF0FFF0FFF1FFF1FFF2FFF2FFF2FFF3FFF3FFF4FFF4FFF5FFF5FFF5FFF6FFF6",
		INIT_70=>X"FFEAFFEBFFEBFFEBFFECFFECFFECFFEDFFEDFFEDFFEEFFEEFFEEFFEFFFEFFFF0",
		INIT_71=>X"FFE7FFE7FFE7FFE7FFE7FFE7FFE8FFE8FFE8FFE8FFE9FFE9FFE9FFE9FFEAFFEA",
		INIT_72=>X"FFE5FFE5FFE5FFE5FFE5FFE5FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6",
		INIT_73=>X"FFE7FFE7FFE7FFE7FFE7FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE5FFE5",
		INIT_74=>X"FFEDFFECFFECFFEBFFEBFFEBFFEAFFEAFFEAFFE9FFE9FFE9FFE8FFE8FFE8FFE8",
		INIT_75=>X"FFF5FFF4FFF4FFF3FFF3FFF2FFF1FFF1FFF0FFF0FFEFFFEFFFEEFFEEFFEDFFED",
		INIT_76=>X"00010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8FFF7FFF6FFF6",
		INIT_77=>X"000F000E000D000C000B000A0009000800070006000600050004000300020001",
		INIT_78=>X"001E001D001C001B001A0019001800170016001500140013001200110010000F",
		INIT_79=>X"002F002E002D002C002B002A002900280027002600250024002200210020001F",
		INIT_7A=>X"0040003F003E003D003C003B0039003800370036003500340033003200310030",
		INIT_7B=>X"004F004E004D004C004B004A0049004900480047004600450044004300420041",
		INIT_7C=>X"005C005C005B005A005900580058005700560055005400530053005200510050",
		INIT_7D=>X"006700660065006500640064006300620062006100610060005F005E005E005D",
		INIT_7E=>X"006D006D006C006C006C006B006B006B006A006A006900690069006800680067",
		INIT_7F=>X"006F006F006F006F006F006F006F006F006F006F006E006E006E006E006E006D",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_01,
		DOPADOP=>dopadop_01,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_02: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000",
		INITP_02=>X"0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFF",
		INITP_03=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000",
		INITP_04=>X"000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_05=>X"FFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000",
		INITP_06=>X"000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_08=>X"FFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000",
		INITP_09=>X"00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0A=>X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000",
		INITP_0B=>X"FFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000",
		INITP_0C=>X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0D=>X"000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000",
		INITP_0F=>X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
		INIT_00=>X"006E006E006E006E006E006F006F006F006F006F006F006F006F006F006F0070",
		INIT_01=>X"00680068006900690069006A006A006B006B006B006C006C006C006D006D006D",
		INIT_02=>X"005E005E005F0060006100610062006200630064006400650065006600670067",
		INIT_03=>X"00510052005300530054005500560057005800580059005A005B005C005C005D",
		INIT_04=>X"004200430044004500460047004800490049004A004B004C004D004E004F0050",
		INIT_05=>X"003100320033003400350036003700380039003B003C003D003E003F00400041",
		INIT_06=>X"002000210022002400250026002700280029002A002B002C002D002E002F0030",
		INIT_07=>X"0010001100120013001400150016001700180019001A001B001C001D001E001F",
		INIT_08=>X"000200030004000500060006000700080009000A000B000C000D000E000F000F",
		INIT_09=>X"FFF6FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFCFFFDFFFDFFFEFFFF000000010001",
		INIT_0A=>X"FFEDFFEEFFEEFFEFFFEFFFF0FFF0FFF1FFF1FFF2FFF3FFF3FFF4FFF4FFF5FFF6",
		INIT_0B=>X"FFE8FFE8FFE8FFE9FFE9FFE9FFEAFFEAFFEAFFEBFFEBFFEBFFECFFECFFEDFFED",
		INIT_0C=>X"FFE5FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE7FFE7FFE7FFE7FFE7FFE8",
		INIT_0D=>X"FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE5FFE5FFE5FFE5FFE5FFE5FFE5",
		INIT_0E=>X"FFEAFFE9FFE9FFE9FFE9FFE8FFE8FFE8FFE8FFE7FFE7FFE7FFE7FFE7FFE7FFE6",
		INIT_0F=>X"FFEFFFEFFFEEFFEEFFEEFFEDFFEDFFEDFFECFFECFFECFFEBFFEBFFEBFFEAFFEA",
		INIT_10=>X"FFF6FFF5FFF5FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF2FFF1FFF1FFF0FFF0FFF0",
		INIT_11=>X"FFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF7FFF7FFF6",
		INIT_12=>X"00040004000300030002000200010001000100000000FFFFFFFFFFFEFFFEFFFD",
		INIT_13=>X"000A000A00090009000900080008000700070007000600060006000500050004",
		INIT_14=>X"000E000E000E000E000D000D000D000D000C000C000C000B000B000B000B000A",
		INIT_15=>X"0011001100110010001000100010001000100010000F000F000F000F000F000E",
		INIT_16=>X"0011001100110011001100110011001100110011001100110011001100110011",
		INIT_17=>X"0010001000100010001000100010001100110011001100110011001100110011",
		INIT_18=>X"000C000D000D000D000D000E000E000E000E000E000F000F000F000F000F0010",
		INIT_19=>X"000800080008000900090009000A000A000A000A000B000B000B000C000C000C",
		INIT_1A=>X"0002000300030003000400040004000500050005000600060006000700070007",
		INIT_1B=>X"FFFDFFFDFFFDFFFEFFFEFFFEFFFFFFFFFFFF0000000000010001000100020002",
		INIT_1C=>X"FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFC",
		INIT_1D=>X"FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_1E=>X"FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3FFF3",
		INIT_1F=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_20=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_21=>X"FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF0",
		INIT_22=>X"FFF7FFF7FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3",
		INIT_23=>X"FFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF7FFF7",
		INIT_24=>X"000200010001000100000000FFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFC",
		INIT_25=>X"0007000700060006000600050005000500040004000400030003000300020002",
		INIT_26=>X"000C000C000B000B000B000A000A000A000A0009000900090008000800080007",
		INIT_27=>X"000F000F000F000F000F000E000E000E000E000E000D000D000D000D000C000C",
		INIT_28=>X"0011001100110011001100110011001100100010001000100010001000100010",
		INIT_29=>X"0011001100110011001100110011001100110011001100110011001100110011",
		INIT_2A=>X"000F000F000F000F000F00100010001000100010001000100011001100110011",
		INIT_2B=>X"000B000B000B000B000C000C000C000D000D000D000D000E000E000E000E000E",
		INIT_2C=>X"0005000500060006000600070007000700080008000900090009000A000A000A",
		INIT_2D=>X"FFFEFFFEFFFFFFFF000000000001000100010002000200030003000400040004",
		INIT_2E=>X"FFF7FFF7FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFD",
		INIT_2F=>X"FFF0FFF0FFF1FFF1FFF2FFF2FFF2FFF3FFF3FFF4FFF4FFF5FFF5FFF5FFF6FFF6",
		INIT_30=>X"FFEAFFEBFFEBFFEBFFECFFECFFECFFEDFFEDFFEDFFEEFFEEFFEEFFEFFFEFFFF0",
		INIT_31=>X"FFE7FFE7FFE7FFE7FFE7FFE7FFE8FFE8FFE8FFE8FFE9FFE9FFE9FFE9FFEAFFEA",
		INIT_32=>X"FFE5FFE5FFE5FFE5FFE5FFE5FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6",
		INIT_33=>X"FFE7FFE7FFE7FFE7FFE7FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE6FFE5FFE5",
		INIT_34=>X"FFEDFFECFFECFFEBFFEBFFEBFFEAFFEAFFEAFFE9FFE9FFE9FFE8FFE8FFE8FFE8",
		INIT_35=>X"FFF5FFF4FFF4FFF3FFF3FFF2FFF1FFF1FFF0FFF0FFEFFFEFFFEEFFEEFFEDFFED",
		INIT_36=>X"00010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8FFF7FFF6FFF6",
		INIT_37=>X"000F000E000D000C000B000A0009000800070006000600050004000300020001",
		INIT_38=>X"001E001D001C001B001A0019001800170016001500140013001200110010000F",
		INIT_39=>X"002F002E002D002C002B002A002900280027002600250024002200210020001F",
		INIT_3A=>X"0040003F003E003D003C003B0039003800370036003500340033003200310030",
		INIT_3B=>X"004F004E004D004C004B004A0049004900480047004600450044004300420041",
		INIT_3C=>X"005C005C005B005A005900580058005700560055005400530053005200510050",
		INIT_3D=>X"006700660065006500640064006300620062006100610060005F005E005E005D",
		INIT_3E=>X"006D006D006C006C006C006B006B006B006A006A006900690069006800680067",
		INIT_3F=>X"006F006F006F006F006F006F006F006F006F006F006E006E006E006E006E006D",
		INIT_40=>X"00A800A900AA00AB00AC00AC00AD00AD00AE00AE00AF00AF00AF00AF00AF00B0",
		INIT_41=>X"00910093009500970098009A009C009D009E00A000A100A300A400A500A600A7",
		INIT_42=>X"006F0071007400760078007B007D007F0081008300850088008A008C008E008F",
		INIT_43=>X"00460049004B004E0051005300560058005B005D0060006300650068006A006C",
		INIT_44=>X"001E0020002300250028002A002D002F0032003400370039003C003F00410044",
		INIT_45=>X"FFFCFFFE00000002000400060008000A000C000E00100012001500170019001C",
		INIT_46=>X"FFE4FFE5FFE7FFE8FFE9FFEAFFECFFEDFFEFFFF0FFF2FFF3FFF5FFF7FFF8FFFA",
		INIT_47=>X"FFD9FFD9FFDAFFDAFFDBFFDBFFDCFFDCFFDDFFDEFFDFFFDFFFE0FFE1FFE2FFE3",
		INIT_48=>X"FFDAFFDAFFD9FFD9FFD9FFD9FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD9FFD9",
		INIT_49=>X"FFE4FFE4FFE3FFE2FFE1FFE0FFE0FFDFFFDEFFDEFFDDFFDCFFDCFFDBFFDBFFDA",
		INIT_4A=>X"FFF4FFF3FFF2FFF1FFF0FFEFFFEEFFEDFFECFFEBFFEAFFE9FFE8FFE7FFE6FFE5",
		INIT_4B=>X"00040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5",
		INIT_4C=>X"001100100010000F000E000E000D000C000B000A000A00090008000700060005",
		INIT_4D=>X"0017001700170017001600160016001500150015001400140013001300120012",
		INIT_4E=>X"0017001700170018001800180018001800180018001800180018001800180018",
		INIT_4F=>X"0010001100110012001200130013001400140015001500150016001600160017",
		INIT_50=>X"000500060007000800080009000A000A000B000C000C000D000E000E000F0010",
		INIT_51=>X"FFFAFFFBFFFBFFFCFFFDFFFEFFFEFFFF00000000000100020003000300040005",
		INIT_52=>X"FFF1FFF2FFF2FFF3FFF3FFF4FFF4FFF5FFF5FFF6FFF6FFF7FFF8FFF8FFF9FFF9",
		INIT_53=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF0FFF1",
		INIT_54=>X"FFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFECFFECFFECFFECFFECFFEDFFED",
		INIT_55=>X"FFF4FFF3FFF3FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFEFFFEFFFEFFFEEFFEEFFEE",
		INIT_56=>X"FFFCFFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF6FFF6FFF5FFF4FFF4",
		INIT_57=>X"00060005000400040003000300020002000100000000FFFFFFFFFFFEFFFDFFFD",
		INIT_58=>X"000D000C000C000C000B000B000A000A000A0009000900080008000700070006",
		INIT_59=>X"001000100010001000100010000F000F000F000F000F000E000E000E000D000D",
		INIT_5A=>X"000F000F000F000F000F00100010001000100010001000100010001000100010",
		INIT_5B=>X"00090009000A000A000B000B000C000C000C000D000D000D000E000E000E000E",
		INIT_5C=>X"0001000100020002000300040004000500050006000600070007000800080009",
		INIT_5D=>X"FFF8FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFEFFFEFFFFFFFF00000000",
		INIT_5E=>X"FFF2FFF2FFF3FFF3FFF3FFF4FFF4FFF4FFF5FFF5FFF6FFF6FFF7FFF7FFF7FFF8",
		INIT_5F=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2",
		INIT_60=>X"FFF1FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_61=>X"FFF7FFF7FFF7FFF6FFF6FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF2FFF2FFF2",
		INIT_62=>X"0000FFFFFFFFFFFEFFFEFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF8FFF8",
		INIT_63=>X"0008000800070007000600060005000500040004000300020002000100010000",
		INIT_64=>X"000E000E000E000D000D000D000C000C000C000B000B000A000A000900090009",
		INIT_65=>X"0010001000100010001000100010001000100010000F000F000F000F000F000E",
		INIT_66=>X"000D000E000E000E000F000F000F000F000F0010001000100010001000100010",
		INIT_67=>X"000700070008000800090009000A000A000A000B000B000C000C000C000D000D",
		INIT_68=>X"FFFDFFFEFFFFFFFF000000000001000200020003000300040004000500060006",
		INIT_69=>X"FFF4FFF5FFF6FFF6FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFCFFFD",
		INIT_6A=>X"FFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF0FFF1FFF1FFF2FFF2FFF3FFF3FFF4FFF4",
		INIT_6B=>X"FFEDFFECFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEEFFEE",
		INIT_6C=>X"FFF0FFF0FFF0FFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFED",
		INIT_6D=>X"FFF9FFF8FFF8FFF7FFF6FFF6FFF5FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF1FFF1",
		INIT_6E=>X"0004000300030002000100000000FFFFFFFEFFFEFFFDFFFCFFFBFFFBFFFAFFF9",
		INIT_6F=>X"000F000E000E000D000C000C000B000A000A0009000800080007000600050005",
		INIT_70=>X"0016001600160015001500150014001400130013001200120011001100100010",
		INIT_71=>X"0018001800180018001800180018001800180018001800180017001700170017",
		INIT_72=>X"0012001300130014001400150015001500160016001600170017001700170018",
		INIT_73=>X"0006000700080009000A000A000B000C000D000E000E000F0010001000110012",
		INIT_74=>X"FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF000000010002000300040005",
		INIT_75=>X"FFE6FFE7FFE8FFE9FFEAFFEBFFECFFEDFFEEFFEFFFF0FFF1FFF2FFF3FFF4FFF5",
		INIT_76=>X"FFDBFFDBFFDCFFDCFFDDFFDEFFDEFFDFFFE0FFE0FFE1FFE2FFE3FFE4FFE4FFE5",
		INIT_77=>X"FFD9FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD9FFD9FFD9FFD9FFDAFFDAFFDA",
		INIT_78=>X"FFE2FFE1FFE0FFDFFFDFFFDEFFDDFFDCFFDCFFDBFFDBFFDAFFDAFFD9FFD9FFD9",
		INIT_79=>X"FFF8FFF7FFF5FFF3FFF2FFF0FFEFFFEDFFECFFEAFFE9FFE8FFE7FFE5FFE4FFE3",
		INIT_7A=>X"00190017001500120010000E000C000A00080006000400020000FFFEFFFCFFFA",
		INIT_7B=>X"0041003F003C0039003700340032002F002D002A0028002500230020001E001C",
		INIT_7C=>X"006A0068006500630060005D005B0058005600530051004E004B004900460044",
		INIT_7D=>X"008E008C008A0088008500830081007F007D007B0078007600740071006F006C",
		INIT_7E=>X"00A600A500A400A300A100A0009E009D009C009A00980097009500930091008F",
		INIT_7F=>X"00AF00AF00AF00AF00AF00AE00AE00AD00AD00AC00AC00AB00AA00A900A800A7",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_02,
		DOPADOP=>dopadop_02,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_03: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000",
		INITP_01=>X"00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_02=>X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000",
		INITP_03=>X"FFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000",
		INITP_04=>X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
		INITP_05=>X"000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000",
		INITP_06=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000",
		INITP_07=>X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
		INITP_08=>X"0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000",
		INITP_09=>X"00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000",
		INITP_0A=>X"00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000",
		INITP_0B=>X"000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000",
		INITP_0C=>X"0000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000",
		INITP_0D=>X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000",
		INITP_0E=>X"00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000",
		INITP_0F=>X"000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000",
		INIT_00=>X"00A800A900AA00AB00AC00AC00AD00AD00AE00AE00AF00AF00AF00AF00AF00B0",
		INIT_01=>X"00910093009500970098009A009C009D009E00A000A100A300A400A500A600A7",
		INIT_02=>X"006F0071007400760078007B007D007F0081008300850088008A008C008E008F",
		INIT_03=>X"00460049004B004E0051005300560058005B005D0060006300650068006A006C",
		INIT_04=>X"001E0020002300250028002A002D002F0032003400370039003C003F00410044",
		INIT_05=>X"FFFCFFFE00000002000400060008000A000C000E00100012001500170019001C",
		INIT_06=>X"FFE4FFE5FFE7FFE8FFE9FFEAFFECFFEDFFEFFFF0FFF2FFF3FFF5FFF7FFF8FFFA",
		INIT_07=>X"FFD9FFD9FFDAFFDAFFDBFFDBFFDCFFDCFFDDFFDEFFDFFFDFFFE0FFE1FFE2FFE3",
		INIT_08=>X"FFDAFFDAFFD9FFD9FFD9FFD9FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD9FFD9",
		INIT_09=>X"FFE4FFE4FFE3FFE2FFE1FFE0FFE0FFDFFFDEFFDEFFDDFFDCFFDCFFDBFFDBFFDA",
		INIT_0A=>X"FFF4FFF3FFF2FFF1FFF0FFEFFFEEFFEDFFECFFEBFFEAFFE9FFE8FFE7FFE6FFE5",
		INIT_0B=>X"00040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5",
		INIT_0C=>X"001100100010000F000E000E000D000C000B000A000A00090008000700060005",
		INIT_0D=>X"0017001700170017001600160016001500150015001400140013001300120012",
		INIT_0E=>X"0017001700170018001800180018001800180018001800180018001800180018",
		INIT_0F=>X"0010001100110012001200130013001400140015001500150016001600160017",
		INIT_10=>X"000500060007000800080009000A000A000B000C000C000D000E000E000F0010",
		INIT_11=>X"FFFAFFFBFFFBFFFCFFFDFFFEFFFEFFFF00000000000100020003000300040005",
		INIT_12=>X"FFF1FFF2FFF2FFF3FFF3FFF4FFF4FFF5FFF5FFF6FFF6FFF7FFF8FFF8FFF9FFF9",
		INIT_13=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF0FFF1",
		INIT_14=>X"FFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFECFFECFFECFFECFFECFFEDFFED",
		INIT_15=>X"FFF4FFF3FFF3FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFEFFFEFFFEFFFEEFFEEFFEE",
		INIT_16=>X"FFFCFFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF6FFF6FFF5FFF4FFF4",
		INIT_17=>X"00060005000400040003000300020002000100000000FFFFFFFFFFFEFFFDFFFD",
		INIT_18=>X"000D000C000C000C000B000B000A000A000A0009000900080008000700070006",
		INIT_19=>X"001000100010001000100010000F000F000F000F000F000E000E000E000D000D",
		INIT_1A=>X"000F000F000F000F000F00100010001000100010001000100010001000100010",
		INIT_1B=>X"00090009000A000A000B000B000C000C000C000D000D000D000E000E000E000E",
		INIT_1C=>X"0001000100020002000300040004000500050006000600070007000800080009",
		INIT_1D=>X"FFF8FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFEFFFEFFFFFFFF00000000",
		INIT_1E=>X"FFF2FFF2FFF3FFF3FFF3FFF4FFF4FFF4FFF5FFF5FFF6FFF6FFF7FFF7FFF7FFF8",
		INIT_1F=>X"FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2",
		INIT_20=>X"FFF1FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_21=>X"FFF7FFF7FFF7FFF6FFF6FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF2FFF2FFF2",
		INIT_22=>X"0000FFFFFFFFFFFEFFFEFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF8FFF8",
		INIT_23=>X"0008000800070007000600060005000500040004000300020002000100010000",
		INIT_24=>X"000E000E000E000D000D000D000C000C000C000B000B000A000A000900090009",
		INIT_25=>X"0010001000100010001000100010001000100010000F000F000F000F000F000E",
		INIT_26=>X"000D000E000E000E000F000F000F000F000F0010001000100010001000100010",
		INIT_27=>X"000700070008000800090009000A000A000A000B000B000C000C000C000D000D",
		INIT_28=>X"FFFDFFFEFFFFFFFF000000000001000200020003000300040004000500060006",
		INIT_29=>X"FFF4FFF5FFF6FFF6FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFCFFFD",
		INIT_2A=>X"FFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF0FFF1FFF1FFF2FFF2FFF3FFF3FFF4FFF4",
		INIT_2B=>X"FFEDFFECFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEEFFEE",
		INIT_2C=>X"FFF0FFF0FFF0FFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFED",
		INIT_2D=>X"FFF9FFF8FFF8FFF7FFF6FFF6FFF5FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF1FFF1",
		INIT_2E=>X"0004000300030002000100000000FFFFFFFEFFFEFFFDFFFCFFFBFFFBFFFAFFF9",
		INIT_2F=>X"000F000E000E000D000C000C000B000A000A0009000800080007000600050005",
		INIT_30=>X"0016001600160015001500150014001400130013001200120011001100100010",
		INIT_31=>X"0018001800180018001800180018001800180018001800180017001700170017",
		INIT_32=>X"0012001300130014001400150015001500160016001600170017001700170018",
		INIT_33=>X"0006000700080009000A000A000B000C000D000E000E000F0010001000110012",
		INIT_34=>X"FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF000000010002000300040005",
		INIT_35=>X"FFE6FFE7FFE8FFE9FFEAFFEBFFECFFEDFFEEFFEFFFF0FFF1FFF2FFF3FFF4FFF5",
		INIT_36=>X"FFDBFFDBFFDCFFDCFFDDFFDEFFDEFFDFFFE0FFE0FFE1FFE2FFE3FFE4FFE4FFE5",
		INIT_37=>X"FFD9FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD9FFD9FFD9FFD9FFDAFFDAFFDA",
		INIT_38=>X"FFE2FFE1FFE0FFDFFFDFFFDEFFDDFFDCFFDCFFDBFFDBFFDAFFDAFFD9FFD9FFD9",
		INIT_39=>X"FFF8FFF7FFF5FFF3FFF2FFF0FFEFFFEDFFECFFEAFFE9FFE8FFE7FFE5FFE4FFE3",
		INIT_3A=>X"00190017001500120010000E000C000A00080006000400020000FFFEFFFCFFFA",
		INIT_3B=>X"0041003F003C0039003700340032002F002D002A0028002500230020001E001C",
		INIT_3C=>X"006A0068006500630060005D005B0058005600530051004E004B004900460044",
		INIT_3D=>X"008E008C008A0088008500830081007F007D007B0078007600740071006F006C",
		INIT_3E=>X"00A600A500A400A300A100A0009E009D009C009A00980097009500930091008F",
		INIT_3F=>X"00AF00AF00AF00AF00AF00AE00AE00AD00AD00AC00AC00AB00AA00A900A800A7",
		INIT_40=>X"00F500F800FB00FE0101010301060108010A010B010C010E010E010F010F0110",
		INIT_41=>X"00A800AE00B300B900BE00C400C900CE00D300D800DC00E100E500E900ED00F1",
		INIT_42=>X"0046004C00520059005F0065006B00710077007E0084008A00900096009C00A2",
		INIT_43=>X"FFF4FFF8FFFC00010005000A000F00140019001E00240029002F0035003B0040",
		INIT_44=>X"FFC8FFCAFFCBFFCDFFCFFFD1FFD3FFD5FFD8FFDBFFDEFFE1FFE4FFE8FFECFFF0",
		INIT_45=>X"FFC9FFC8FFC7FFC6FFC5FFC5FFC4FFC4FFC4FFC4FFC4FFC4FFC5FFC5FFC6FFC7",
		INIT_46=>X"FFE9FFE6FFE4FFE2FFDFFFDDFFDBFFD9FFD7FFD5FFD3FFD1FFCFFFCEFFCCFFCB",
		INIT_47=>X"000E000C000A0007000500030001FFFEFFFCFFFAFFF7FFF5FFF2FFF0FFEEFFEB",
		INIT_48=>X"0022002200210020001F001E001D001C001B0019001800160015001300110010",
		INIT_49=>X"001E001F00200021002200220023002300230024002400240024002300230023",
		INIT_4A=>X"0009000A000C000D000F0011001200130015001600180019001A001B001C001D",
		INIT_4B=>X"FFF1FFF2FFF3FFF5FFF6FFF7FFF9FFFAFFFCFFFDFFFF00010002000400050007",
		INIT_4C=>X"FFE5FFE5FFE6FFE6FFE6FFE7FFE7FFE8FFE9FFEAFFEAFFEBFFECFFEDFFEEFFF0",
		INIT_4D=>X"FFEBFFEAFFEAFFE9FFE8FFE7FFE7FFE6FFE6FFE6FFE5FFE5FFE5FFE5FFE5FFE5",
		INIT_4E=>X"FFFDFFFCFFFBFFF9FFF8FFF7FFF6FFF4FFF3FFF2FFF1FFF0FFEFFFEEFFEDFFEC",
		INIT_4F=>X"000F000E000D000C000B000A000900080007000600040003000200010000FFFE",
		INIT_50=>X"0015001500150015001500150014001400140013001300120012001100100010",
		INIT_51=>X"000D000E000F0010001100110012001200130013001400140014001500150015",
		INIT_52=>X"FFFEFFFF0000000100020003000400050006000700080009000A000B000C000D",
		INIT_53=>X"FFF0FFF1FFF1FFF2FFF3FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFD",
		INIT_54=>X"FFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEFFFEFFFF0",
		INIT_55=>X"FFF6FFF5FFF5FFF4FFF3FFF2FFF2FFF1FFF0FFF0FFEFFFEFFFEEFFEEFFEEFFED",
		INIT_56=>X"000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF7",
		INIT_57=>X"000F000F000E000E000D000D000C000C000B000A000900090008000700060005",
		INIT_58=>X"000F001000100010001000100011001100110011001100100010001000100010",
		INIT_59=>X"000500060007000800080009000A000B000B000C000C000D000D000E000E000F",
		INIT_5A=>X"FFF8FFF9FFF9FFFAFFFBFFFCFFFDFFFDFFFEFFFF000000010002000300040004",
		INIT_5B=>X"FFF0FFF0FFF0FFF0FFF1FFF1FFF2FFF2FFF3FFF3FFF4FFF4FFF5FFF6FFF6FFF7",
		INIT_5C=>X"FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEFFFEFFFF0",
		INIT_5D=>X"FFFDFFFCFFFBFFFBFFFAFFF9FFF8FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF3FFF3",
		INIT_5E=>X"000A0009000800080007000600050005000400030002000100000000FFFFFFFE",
		INIT_5F=>X"000F000F000F000F000F000F000E000E000E000D000D000C000C000B000B000A",
		INIT_60=>X"000B000B000C000C000D000D000E000E000E000F000F000F000F000F000F0010",
		INIT_61=>X"FFFF0000000000010002000300040005000500060007000800080009000A000A",
		INIT_62=>X"FFF3FFF4FFF4FFF5FFF5FFF6FFF7FFF8FFF8FFF9FFFAFFFBFFFBFFFCFFFDFFFE",
		INIT_63=>X"FFEFFFEFFFEFFFEFFFEFFFEFFFEFFFF0FFF0FFF0FFF0FFF1FFF1FFF2FFF2FFF3",
		INIT_64=>X"FFF6FFF6FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFF0FFF0",
		INIT_65=>X"00040003000200010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF7",
		INIT_66=>X"000E000E000D000D000C000C000B000B000A0009000800080007000600050004",
		INIT_67=>X"00100010001000100011001100110011001100100010001000100010000F000F",
		INIT_68=>X"00060007000800090009000A000B000C000C000D000D000E000E000F000F0010",
		INIT_69=>X"FFF8FFF9FFFAFFFAFFFBFFFCFFFDFFFEFFFF0000000100020003000400050005",
		INIT_6A=>X"FFEEFFEEFFEEFFEFFFEFFFF0FFF0FFF1FFF2FFF2FFF3FFF4FFF5FFF5FFF6FFF7",
		INIT_6B=>X"FFEFFFEFFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFED",
		INIT_6C=>X"FFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF3FFF3FFF2FFF1FFF1FFF0FFF0",
		INIT_6D=>X"000C000B000A0009000800070006000500040003000200010000FFFFFFFEFFFD",
		INIT_6E=>X"001500150014001400140013001300120012001100110010000F000E000D000D",
		INIT_6F=>X"0010001100120012001300130014001400140015001500150015001500150015",
		INIT_70=>X"000000010002000300040006000700080009000A000B000C000D000E000F0010",
		INIT_71=>X"FFEDFFEEFFEFFFF0FFF1FFF2FFF3FFF4FFF6FFF7FFF8FFF9FFFBFFFCFFFDFFFE",
		INIT_72=>X"FFE5FFE5FFE5FFE5FFE5FFE6FFE6FFE6FFE7FFE7FFE8FFE9FFEAFFEAFFEBFFEC",
		INIT_73=>X"FFEEFFEDFFECFFEBFFEAFFEAFFE9FFE8FFE7FFE7FFE6FFE6FFE6FFE5FFE5FFE5",
		INIT_74=>X"0005000400020001FFFFFFFDFFFCFFFAFFF9FFF7FFF6FFF5FFF3FFF2FFF1FFF0",
		INIT_75=>X"001C001B001A0019001800160015001300120011000F000D000C000A00090007",
		INIT_76=>X"0023002300240024002400240023002300230022002200210020001F001E001D",
		INIT_77=>X"001100130015001600180019001B001C001D001E001F00200021002200220023",
		INIT_78=>X"FFEEFFF0FFF2FFF5FFF7FFFAFFFCFFFE0001000300050007000A000C000E0010",
		INIT_79=>X"FFCCFFCEFFCFFFD1FFD3FFD5FFD7FFD9FFDBFFDDFFDFFFE2FFE4FFE6FFE9FFEB",
		INIT_7A=>X"FFC6FFC5FFC5FFC4FFC4FFC4FFC4FFC4FFC4FFC5FFC5FFC6FFC7FFC8FFC9FFCB",
		INIT_7B=>X"FFECFFE8FFE4FFE1FFDEFFDBFFD8FFD5FFD3FFD1FFCFFFCDFFCBFFCAFFC8FFC7",
		INIT_7C=>X"003B0035002F00290024001E00190014000F000A00050001FFFCFFF8FFF4FFF0",
		INIT_7D=>X"009C00960090008A0084007E00770071006B0065005F00590052004C00460040",
		INIT_7E=>X"00ED00E900E500E100DC00D800D300CE00C900C400BE00B900B300AE00A800A2",
		INIT_7F=>X"010F010F010E010E010C010B010A010801060103010100FE00FB00F800F500F1",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_03,
		DOPADOP=>dopadop_03,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_04: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000",
		INITP_01=>X"00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000",
		INITP_02=>X"00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000",
		INITP_03=>X"000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000",
		INITP_04=>X"0000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000",
		INITP_05=>X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000",
		INITP_06=>X"00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000",
		INITP_07=>X"000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000",
		INITP_08=>X"FFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000",
		INITP_09=>X"00000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFF",
		INITP_0A=>X"FFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC000000000000000",
		INITP_0B=>X"0000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFF",
		INITP_0C=>X"FFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC0000000000",
		INITP_0D=>X"000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFF",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000",
		INITP_0F=>X"00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFF",
		INIT_00=>X"00F500F800FB00FE0101010301060108010A010B010C010E010E010F010F0110",
		INIT_01=>X"00A800AE00B300B900BE00C400C900CE00D300D800DC00E100E500E900ED00F1",
		INIT_02=>X"0046004C00520059005F0065006B00710077007E0084008A00900096009C00A2",
		INIT_03=>X"FFF4FFF8FFFC00010005000A000F00140019001E00240029002F0035003B0040",
		INIT_04=>X"FFC8FFCAFFCBFFCDFFCFFFD1FFD3FFD5FFD8FFDBFFDEFFE1FFE4FFE8FFECFFF0",
		INIT_05=>X"FFC9FFC8FFC7FFC6FFC5FFC5FFC4FFC4FFC4FFC4FFC4FFC4FFC5FFC5FFC6FFC7",
		INIT_06=>X"FFE9FFE6FFE4FFE2FFDFFFDDFFDBFFD9FFD7FFD5FFD3FFD1FFCFFFCEFFCCFFCB",
		INIT_07=>X"000E000C000A0007000500030001FFFEFFFCFFFAFFF7FFF5FFF2FFF0FFEEFFEB",
		INIT_08=>X"0022002200210020001F001E001D001C001B0019001800160015001300110010",
		INIT_09=>X"001E001F00200021002200220023002300230024002400240024002300230023",
		INIT_0A=>X"0009000A000C000D000F0011001200130015001600180019001A001B001C001D",
		INIT_0B=>X"FFF1FFF2FFF3FFF5FFF6FFF7FFF9FFFAFFFCFFFDFFFF00010002000400050007",
		INIT_0C=>X"FFE5FFE5FFE6FFE6FFE6FFE7FFE7FFE8FFE9FFEAFFEAFFEBFFECFFEDFFEEFFF0",
		INIT_0D=>X"FFEBFFEAFFEAFFE9FFE8FFE7FFE7FFE6FFE6FFE6FFE5FFE5FFE5FFE5FFE5FFE5",
		INIT_0E=>X"FFFDFFFCFFFBFFF9FFF8FFF7FFF6FFF4FFF3FFF2FFF1FFF0FFEFFFEEFFEDFFEC",
		INIT_0F=>X"000F000E000D000C000B000A000900080007000600040003000200010000FFFE",
		INIT_10=>X"0015001500150015001500150014001400140013001300120012001100100010",
		INIT_11=>X"000D000E000F0010001100110012001200130013001400140014001500150015",
		INIT_12=>X"FFFEFFFF0000000100020003000400050006000700080009000A000B000C000D",
		INIT_13=>X"FFF0FFF1FFF1FFF2FFF3FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFD",
		INIT_14=>X"FFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEFFFEFFFF0",
		INIT_15=>X"FFF6FFF5FFF5FFF4FFF3FFF2FFF2FFF1FFF0FFF0FFEFFFEFFFEEFFEEFFEEFFED",
		INIT_16=>X"000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF7",
		INIT_17=>X"000F000F000E000E000D000D000C000C000B000A000900090008000700060005",
		INIT_18=>X"000F001000100010001000100011001100110011001100100010001000100010",
		INIT_19=>X"000500060007000800080009000A000B000B000C000C000D000D000E000E000F",
		INIT_1A=>X"FFF8FFF9FFF9FFFAFFFBFFFCFFFDFFFDFFFEFFFF000000010002000300040004",
		INIT_1B=>X"FFF0FFF0FFF0FFF0FFF1FFF1FFF2FFF2FFF3FFF3FFF4FFF4FFF5FFF6FFF6FFF7",
		INIT_1C=>X"FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEFFFEFFFF0",
		INIT_1D=>X"FFFDFFFCFFFBFFFBFFFAFFF9FFF8FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF3FFF3",
		INIT_1E=>X"000A0009000800080007000600050005000400030002000100000000FFFFFFFE",
		INIT_1F=>X"000F000F000F000F000F000F000E000E000E000D000D000C000C000B000B000A",
		INIT_20=>X"000B000B000C000C000D000D000E000E000E000F000F000F000F000F000F0010",
		INIT_21=>X"FFFF0000000000010002000300040005000500060007000800080009000A000A",
		INIT_22=>X"FFF3FFF4FFF4FFF5FFF5FFF6FFF7FFF8FFF8FFF9FFFAFFFBFFFBFFFCFFFDFFFE",
		INIT_23=>X"FFEFFFEFFFEFFFEFFFEFFFEFFFEFFFF0FFF0FFF0FFF0FFF1FFF1FFF2FFF2FFF3",
		INIT_24=>X"FFF6FFF6FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFF0FFF0",
		INIT_25=>X"00040003000200010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF7",
		INIT_26=>X"000E000E000D000D000C000C000B000B000A0009000800080007000600050004",
		INIT_27=>X"00100010001000100011001100110011001100100010001000100010000F000F",
		INIT_28=>X"00060007000800090009000A000B000C000C000D000D000E000E000F000F0010",
		INIT_29=>X"FFF8FFF9FFFAFFFAFFFBFFFCFFFDFFFEFFFF0000000100020003000400050005",
		INIT_2A=>X"FFEEFFEEFFEEFFEFFFEFFFF0FFF0FFF1FFF2FFF2FFF3FFF4FFF5FFF5FFF6FFF7",
		INIT_2B=>X"FFEFFFEFFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFED",
		INIT_2C=>X"FFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF3FFF3FFF2FFF1FFF1FFF0FFF0",
		INIT_2D=>X"000C000B000A0009000800070006000500040003000200010000FFFFFFFEFFFD",
		INIT_2E=>X"001500150014001400140013001300120012001100110010000F000E000D000D",
		INIT_2F=>X"0010001100120012001300130014001400140015001500150015001500150015",
		INIT_30=>X"000000010002000300040006000700080009000A000B000C000D000E000F0010",
		INIT_31=>X"FFEDFFEEFFEFFFF0FFF1FFF2FFF3FFF4FFF6FFF7FFF8FFF9FFFBFFFCFFFDFFFE",
		INIT_32=>X"FFE5FFE5FFE5FFE5FFE5FFE6FFE6FFE6FFE7FFE7FFE8FFE9FFEAFFEAFFEBFFEC",
		INIT_33=>X"FFEEFFEDFFECFFEBFFEAFFEAFFE9FFE8FFE7FFE7FFE6FFE6FFE6FFE5FFE5FFE5",
		INIT_34=>X"0005000400020001FFFFFFFDFFFCFFFAFFF9FFF7FFF6FFF5FFF3FFF2FFF1FFF0",
		INIT_35=>X"001C001B001A0019001800160015001300120011000F000D000C000A00090007",
		INIT_36=>X"0023002300240024002400240023002300230022002200210020001F001E001D",
		INIT_37=>X"001100130015001600180019001B001C001D001E001F00200021002200220023",
		INIT_38=>X"FFEEFFF0FFF2FFF5FFF7FFFAFFFCFFFE0001000300050007000A000C000E0010",
		INIT_39=>X"FFCCFFCEFFCFFFD1FFD3FFD5FFD7FFD9FFDBFFDDFFDFFFE2FFE4FFE6FFE9FFEB",
		INIT_3A=>X"FFC6FFC5FFC5FFC4FFC4FFC4FFC4FFC4FFC4FFC5FFC5FFC6FFC7FFC8FFC9FFCB",
		INIT_3B=>X"FFECFFE8FFE4FFE1FFDEFFDBFFD8FFD5FFD3FFD1FFCFFFCDFFCBFFCAFFC8FFC7",
		INIT_3C=>X"003B0035002F00290024001E00190014000F000A00050001FFFCFFF8FFF4FFF0",
		INIT_3D=>X"009C00960090008A0084007E00770071006B0065005F00590052004C00460040",
		INIT_3E=>X"00ED00E900E500E100DC00D800D300CE00C900C400BE00B900B300AE00A800A2",
		INIT_3F=>X"010F010F010E010E010C010B010A010801060103010100FE00FB00F800F500F1",
		INIT_40=>X"013D0147015101590162016901710177017D018201860189018C018E018F0190",
		INIT_41=>X"00740081008E009C00A900B700C400D100DE00EB00F801040110011C01280133",
		INIT_42=>X"FFCEFFD5FFDCFFE4FFEDFFF6FFFF00090014001E002A00350041004E005A0067",
		INIT_43=>X"FFADFFABFFAAFFA9FFA8FFA8FFA9FFAAFFACFFAEFFB1FFB4FFB8FFBDFFC2FFC7",
		INIT_44=>X"FFF1FFECFFE6FFE1FFDCFFD7FFD2FFCDFFC8FFC4FFC0FFBCFFB8FFB5FFB2FFAF",
		INIT_45=>X"002E002C002A002800250022001E001A00170012000E000900050000FFFBFFF6",
		INIT_46=>X"00250028002A002C002E00300031003200330033003400340033003200310030",
		INIT_47=>X"FFF2FFF5FFF9FFFCFFFF000200060009000D001000130017001A001D00200023",
		INIT_48=>X"FFDAFFDAFFDAFFDAFFDBFFDCFFDDFFDEFFE0FFE1FFE3FFE5FFE8FFEAFFEDFFF0",
		INIT_49=>X"FFF3FFF1FFEEFFECFFEAFFE7FFE5FFE3FFE2FFE0FFDFFFDDFFDCFFDBFFDBFFDA",
		INIT_4A=>X"00170016001400120010000E000C000A0007000500020000FFFDFFFBFFF8FFF6",
		INIT_4B=>X"0019001A001B001C001C001D001D001D001D001D001D001C001C001B001A0018",
		INIT_4C=>X"FFFBFFFDFFFF0001000300050007000A000C000D000F00110013001500160017",
		INIT_4D=>X"FFE7FFE7FFE7FFE8FFE9FFEAFFEBFFECFFEDFFEFFFF0FFF2FFF3FFF5FFF7FFF9",
		INIT_4E=>X"FFF4FFF2FFF1FFEFFFEEFFECFFEBFFEAFFE9FFE8FFE8FFE7FFE7FFE7FFE6FFE6",
		INIT_4F=>X"000E000D000C000A000800070005000300020000FFFEFFFCFFFBFFF9FFF7FFF5",
		INIT_50=>X"0014001400150015001500150015001500150015001400130013001200110010",
		INIT_51=>X"FFFF000100020004000500070008000A000B000D000E000F0010001100120013",
		INIT_52=>X"FFEDFFEDFFEEFFEEFFEFFFF0FFF1FFF2FFF3FFF5FFF6FFF7FFF9FFFAFFFCFFFD",
		INIT_53=>X"FFF4FFF2FFF1FFF0FFEFFFEFFFEEFFEDFFEDFFECFFECFFECFFECFFECFFECFFEC",
		INIT_54=>X"00090008000700060004000300010000FFFFFFFDFFFCFFFAFFF9FFF7FFF6FFF5",
		INIT_55=>X"0011001200120012001200120011001100100010000F000F000E000D000C000B",
		INIT_56=>X"0002000300040006000700080009000B000C000D000E000E000F001000100011",
		INIT_57=>X"FFF0FFF1FFF1FFF2FFF3FFF4FFF5FFF6FFF7FFF8FFFAFFFBFFFCFFFEFFFF0000",
		INIT_58=>X"FFF3FFF2FFF1FFF1FFF0FFF0FFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEFFFEFFFF0",
		INIT_59=>X"000600050004000300010000FFFFFFFDFFFCFFFBFFFAFFF8FFF7FFF6FFF5FFF4",
		INIT_5A=>X"00100010001000100010000F000F000E000E000D000C000B000B000A00080007",
		INIT_5B=>X"000400050006000700080009000A000B000C000D000E000E000F000F00100010",
		INIT_5C=>X"FFF2FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFEFFFF000000010003",
		INIT_5D=>X"FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFEFFFEFFFEFFFF0FFF0FFF0FFF1FFF1FFF2",
		INIT_5E=>X"0004000300010000FFFFFFFEFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF3",
		INIT_5F=>X"000F000F000F000F000E000E000D000D000C000B000A00090008000700060005",
		INIT_60=>X"0006000700080009000A000B000C000D000D000E000E000F000F000F000F0010",
		INIT_61=>X"FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFEFFFF00000001000300040005",
		INIT_62=>X"FFF1FFF1FFF0FFF0FFF0FFEFFFEFFFEFFFF0FFF0FFF0FFF1FFF1FFF2FFF2FFF3",
		INIT_63=>X"00010000FFFFFFFEFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF3FFF2FFF2",
		INIT_64=>X"0010000F000F000E000E000D000C000B000A0009000800070006000500040003",
		INIT_65=>X"0008000A000B000B000C000D000E000E000F000F001000100010001000100010",
		INIT_66=>X"FFF5FFF6FFF7FFF8FFFAFFFBFFFCFFFDFFFF0000000100030004000500060007",
		INIT_67=>X"FFEFFFEFFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF1FFF1FFF2FFF3FFF4",
		INIT_68=>X"FFFFFFFEFFFCFFFBFFFAFFF8FFF7FFF6FFF5FFF4FFF3FFF2FFF1FFF1FFF0FFF0",
		INIT_69=>X"00100010000F000E000E000D000C000B00090008000700060004000300020000",
		INIT_6A=>X"000C000D000E000F000F00100010001100110012001200120012001200110011",
		INIT_6B=>X"FFF6FFF7FFF9FFFAFFFCFFFDFFFF00000001000300040006000700080009000B",
		INIT_6C=>X"FFECFFECFFECFFECFFECFFECFFEDFFEDFFEEFFEFFFEFFFF0FFF1FFF2FFF4FFF5",
		INIT_6D=>X"FFFCFFFAFFF9FFF7FFF6FFF5FFF3FFF2FFF1FFF0FFEFFFEEFFEEFFEDFFEDFFEC",
		INIT_6E=>X"001200110010000F000E000D000B000A000800070005000400020001FFFFFFFD",
		INIT_6F=>X"0011001200130013001400150015001500150015001500150015001400140013",
		INIT_70=>X"FFF7FFF9FFFBFFFCFFFE000000020003000500070008000A000C000D000E0010",
		INIT_71=>X"FFE6FFE7FFE7FFE7FFE8FFE8FFE9FFEAFFEBFFECFFEEFFEFFFF1FFF2FFF4FFF5",
		INIT_72=>X"FFF7FFF5FFF3FFF2FFF0FFEFFFEDFFECFFEBFFEAFFE9FFE8FFE7FFE7FFE7FFE6",
		INIT_73=>X"0016001500130011000F000D000C000A0007000500030001FFFFFFFDFFFBFFF9",
		INIT_74=>X"001A001B001C001C001D001D001D001D001D001D001C001C001B001A00190017",
		INIT_75=>X"FFF8FFFBFFFD0000000200050007000A000C000E001000120014001600170018",
		INIT_76=>X"FFDBFFDBFFDCFFDDFFDFFFE0FFE2FFE3FFE5FFE7FFEAFFECFFEEFFF1FFF3FFF6",
		INIT_77=>X"FFEDFFEAFFE8FFE5FFE3FFE1FFE0FFDEFFDDFFDCFFDBFFDAFFDAFFDAFFDAFFDA",
		INIT_78=>X"0020001D001A001700130010000D000900060002FFFFFFFCFFF9FFF5FFF2FFF0",
		INIT_79=>X"0031003200330034003400330033003200310030002E002C002A002800250023",
		INIT_7A=>X"FFFB000000050009000E00120017001A001E002200250028002A002C002E0030",
		INIT_7B=>X"FFB2FFB5FFB8FFBCFFC0FFC4FFC8FFCDFFD2FFD7FFDCFFE1FFE6FFECFFF1FFF6",
		INIT_7C=>X"FFC2FFBDFFB8FFB4FFB1FFAEFFACFFAAFFA9FFA8FFA8FFA9FFAAFFABFFADFFAF",
		INIT_7D=>X"005A004E00410035002A001E00140009FFFFFFF6FFEDFFE4FFDCFFD5FFCEFFC7",
		INIT_7E=>X"0128011C0110010400F800EB00DE00D100C400B700A9009C008E008100740067",
		INIT_7F=>X"018F018E018C018901860182017D0177017101690162015901510147013D0133",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_04,
		DOPADOP=>dopadop_04,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_05: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000",
		INITP_01=>X"00000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFF",
		INITP_02=>X"FFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC000000000000000",
		INITP_03=>X"0000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFF",
		INITP_04=>X"FFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC0000000000",
		INITP_05=>X"000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFF",
		INITP_06=>X"FFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000",
		INITP_07=>X"00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFF",
		INITP_08=>X"00000FFFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF000000000000000",
		INITP_09=>X"00000000003FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFC000000000",
		INITP_0A=>X"FC00000000000000FFFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF0000",
		INITP_0B=>X"FFFFFFF000000000000003FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFF",
		INITP_0C=>X"FFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFF000000000000003FFFFFFF",
		INITP_0D=>X"0003FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFFC00000000000000FF",
		INITP_0E=>X"000000000FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFF00000000000",
		INITP_0F=>X"000000000000003FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFFC00000",
		INIT_00=>X"013D0147015101590162016901710177017D018201860189018C018E018F0190",
		INIT_01=>X"00740081008E009C00A900B700C400D100DE00EB00F801040110011C01280133",
		INIT_02=>X"FFCEFFD5FFDCFFE4FFEDFFF6FFFF00090014001E002A00350041004E005A0067",
		INIT_03=>X"FFADFFABFFAAFFA9FFA8FFA8FFA9FFAAFFACFFAEFFB1FFB4FFB8FFBDFFC2FFC7",
		INIT_04=>X"FFF1FFECFFE6FFE1FFDCFFD7FFD2FFCDFFC8FFC4FFC0FFBCFFB8FFB5FFB2FFAF",
		INIT_05=>X"002E002C002A002800250022001E001A00170012000E000900050000FFFBFFF6",
		INIT_06=>X"00250028002A002C002E00300031003200330033003400340033003200310030",
		INIT_07=>X"FFF2FFF5FFF9FFFCFFFF000200060009000D001000130017001A001D00200023",
		INIT_08=>X"FFDAFFDAFFDAFFDAFFDBFFDCFFDDFFDEFFE0FFE1FFE3FFE5FFE8FFEAFFEDFFF0",
		INIT_09=>X"FFF3FFF1FFEEFFECFFEAFFE7FFE5FFE3FFE2FFE0FFDFFFDDFFDCFFDBFFDBFFDA",
		INIT_0A=>X"00170016001400120010000E000C000A0007000500020000FFFDFFFBFFF8FFF6",
		INIT_0B=>X"0019001A001B001C001C001D001D001D001D001D001D001C001C001B001A0018",
		INIT_0C=>X"FFFBFFFDFFFF0001000300050007000A000C000D000F00110013001500160017",
		INIT_0D=>X"FFE7FFE7FFE7FFE8FFE9FFEAFFEBFFECFFEDFFEFFFF0FFF2FFF3FFF5FFF7FFF9",
		INIT_0E=>X"FFF4FFF2FFF1FFEFFFEEFFECFFEBFFEAFFE9FFE8FFE8FFE7FFE7FFE7FFE6FFE6",
		INIT_0F=>X"000E000D000C000A000800070005000300020000FFFEFFFCFFFBFFF9FFF7FFF5",
		INIT_10=>X"0014001400150015001500150015001500150015001400130013001200110010",
		INIT_11=>X"FFFF000100020004000500070008000A000B000D000E000F0010001100120013",
		INIT_12=>X"FFEDFFEDFFEEFFEEFFEFFFF0FFF1FFF2FFF3FFF5FFF6FFF7FFF9FFFAFFFCFFFD",
		INIT_13=>X"FFF4FFF2FFF1FFF0FFEFFFEFFFEEFFEDFFEDFFECFFECFFECFFECFFECFFECFFEC",
		INIT_14=>X"00090008000700060004000300010000FFFFFFFDFFFCFFFAFFF9FFF7FFF6FFF5",
		INIT_15=>X"0011001200120012001200120011001100100010000F000F000E000D000C000B",
		INIT_16=>X"0002000300040006000700080009000B000C000D000E000E000F001000100011",
		INIT_17=>X"FFF0FFF1FFF1FFF2FFF3FFF4FFF5FFF6FFF7FFF8FFFAFFFBFFFCFFFEFFFF0000",
		INIT_18=>X"FFF3FFF2FFF1FFF1FFF0FFF0FFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEFFFEFFFF0",
		INIT_19=>X"000600050004000300010000FFFFFFFDFFFCFFFBFFFAFFF8FFF7FFF6FFF5FFF4",
		INIT_1A=>X"00100010001000100010000F000F000E000E000D000C000B000B000A00080007",
		INIT_1B=>X"000400050006000700080009000A000B000C000D000E000E000F000F00100010",
		INIT_1C=>X"FFF2FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFEFFFF000000010003",
		INIT_1D=>X"FFF2FFF2FFF1FFF1FFF0FFF0FFF0FFEFFFEFFFEFFFF0FFF0FFF0FFF1FFF1FFF2",
		INIT_1E=>X"0004000300010000FFFFFFFEFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF3",
		INIT_1F=>X"000F000F000F000F000E000E000D000D000C000B000A00090008000700060005",
		INIT_20=>X"0006000700080009000A000B000C000D000D000E000E000F000F000F000F0010",
		INIT_21=>X"FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFEFFFF00000001000300040005",
		INIT_22=>X"FFF1FFF1FFF0FFF0FFF0FFEFFFEFFFEFFFF0FFF0FFF0FFF1FFF1FFF2FFF2FFF3",
		INIT_23=>X"00010000FFFFFFFEFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF3FFF2FFF2",
		INIT_24=>X"0010000F000F000E000E000D000C000B000A0009000800070006000500040003",
		INIT_25=>X"0008000A000B000B000C000D000E000E000F000F001000100010001000100010",
		INIT_26=>X"FFF5FFF6FFF7FFF8FFFAFFFBFFFCFFFDFFFF0000000100030004000500060007",
		INIT_27=>X"FFEFFFEFFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFF0FFF0FFF1FFF1FFF2FFF3FFF4",
		INIT_28=>X"FFFFFFFEFFFCFFFBFFFAFFF8FFF7FFF6FFF5FFF4FFF3FFF2FFF1FFF1FFF0FFF0",
		INIT_29=>X"00100010000F000E000E000D000C000B00090008000700060004000300020000",
		INIT_2A=>X"000C000D000E000F000F00100010001100110012001200120012001200110011",
		INIT_2B=>X"FFF6FFF7FFF9FFFAFFFCFFFDFFFF00000001000300040006000700080009000B",
		INIT_2C=>X"FFECFFECFFECFFECFFECFFECFFEDFFEDFFEEFFEFFFEFFFF0FFF1FFF2FFF4FFF5",
		INIT_2D=>X"FFFCFFFAFFF9FFF7FFF6FFF5FFF3FFF2FFF1FFF0FFEFFFEEFFEEFFEDFFEDFFEC",
		INIT_2E=>X"001200110010000F000E000D000B000A000800070005000400020001FFFFFFFD",
		INIT_2F=>X"0011001200130013001400150015001500150015001500150015001400140013",
		INIT_30=>X"FFF7FFF9FFFBFFFCFFFE000000020003000500070008000A000C000D000E0010",
		INIT_31=>X"FFE6FFE7FFE7FFE7FFE8FFE8FFE9FFEAFFEBFFECFFEEFFEFFFF1FFF2FFF4FFF5",
		INIT_32=>X"FFF7FFF5FFF3FFF2FFF0FFEFFFEDFFECFFEBFFEAFFE9FFE8FFE7FFE7FFE7FFE6",
		INIT_33=>X"0016001500130011000F000D000C000A0007000500030001FFFFFFFDFFFBFFF9",
		INIT_34=>X"001A001B001C001C001D001D001D001D001D001D001C001C001B001A00190017",
		INIT_35=>X"FFF8FFFBFFFD0000000200050007000A000C000E001000120014001600170018",
		INIT_36=>X"FFDBFFDBFFDCFFDDFFDFFFE0FFE2FFE3FFE5FFE7FFEAFFECFFEEFFF1FFF3FFF6",
		INIT_37=>X"FFEDFFEAFFE8FFE5FFE3FFE1FFE0FFDEFFDDFFDCFFDBFFDAFFDAFFDAFFDAFFDA",
		INIT_38=>X"0020001D001A001700130010000D000900060002FFFFFFFCFFF9FFF5FFF2FFF0",
		INIT_39=>X"0031003200330034003400330033003200310030002E002C002A002800250023",
		INIT_3A=>X"FFFB000000050009000E00120017001A001E002200250028002A002C002E0030",
		INIT_3B=>X"FFB2FFB5FFB8FFBCFFC0FFC4FFC8FFCDFFD2FFD7FFDCFFE1FFE6FFECFFF1FFF6",
		INIT_3C=>X"FFC2FFBDFFB8FFB4FFB1FFAEFFACFFAAFFA9FFA8FFA8FFA9FFAAFFABFFADFFAF",
		INIT_3D=>X"005A004E00410035002A001E00140009FFFFFFF6FFEDFFE4FFDCFFD5FFCEFFC7",
		INIT_3E=>X"0128011C0110010400F800EB00DE00D100C400B700A9009C008E008100740067",
		INIT_3F=>X"018F018E018C018901860182017D0177017101690162015901510147013D0133",
		INIT_40=>X"015B0173018B01A101B601CA01DC01ED01FC020A0215021E0226022B022E0230",
		INIT_41=>X"FFE0FFF200040019002E0044005C0074008D00A600C000DA00F4010F01290142",
		INIT_42=>X"FF96FF91FF8CFF89FF86FF86FF86FF88FF8BFF91FF97FF9FFFA9FFB5FFC2FFD0",
		INIT_43=>X"0026001E0016000D0004FFFBFFF1FFE7FFDCFFD2FFC8FFBFFFB5FFADFFA4FF9D",
		INIT_44=>X"0035003A003E004200440046004800480048004600440041003D00390033002D",
		INIT_45=>X"FFD8FFDDFFE1FFE6FFECFFF2FFF8FFFE0005000B00120018001F0025002B0030",
		INIT_46=>X"FFE3FFDEFFDAFFD7FFD4FFD1FFCFFFCDFFCCFFCCFFCCFFCCFFCEFFCFFFD2FFD5",
		INIT_47=>X"002400220020001D001900160012000D00090004FFFFFFFAFFF5FFF1FFECFFE7",
		INIT_48=>X"000D001000140018001B001E0020002300250026002700280028002800270026",
		INIT_49=>X"FFDEFFDFFFE0FFE1FFE3FFE6FFE8FFEBFFEEFFF2FFF5FFF9FFFD000100050009",
		INIT_4A=>X"FFFEFFFAFFF7FFF4FFF1FFEDFFEBFFE8FFE6FFE3FFE2FFE0FFDFFFDEFFDEFFDE",
		INIT_4B=>X"001C001D001C001C001B001A00190017001500130010000E000B000800040001",
		INIT_4C=>X"FFF9FFFCFFFF000200050008000A000D00100012001400160018001A001B001C",
		INIT_4D=>X"FFE8FFE7FFE6FFE6FFE6FFE6FFE6FFE7FFE8FFEAFFEBFFEDFFEFFFF1FFF4FFF6",
		INIT_4E=>X"000C0009000700050002FFFFFFFDFFFAFFF8FFF5FFF3FFF0FFEEFFECFFEBFFE9",
		INIT_4F=>X"001100130014001500160016001700170016001600150014001300110010000E",
		INIT_50=>X"FFF0FFF1FFF3FFF5FFF7FFF9FFFCFFFE0000000300050007000A000C000E0010",
		INIT_51=>X"FFF4FFF2FFF0FFEFFFEEFFECFFECFFEBFFEAFFEAFFEAFFEBFFEBFFECFFEDFFEE",
		INIT_52=>X"00110010000F000E000C000B00090007000500030000FFFEFFFCFFFAFFF8FFF6",
		INIT_53=>X"000500070009000B000D000E000F001100120012001300130013001300130012",
		INIT_54=>X"FFEDFFEDFFEEFFEFFFF0FFF1FFF2FFF4FFF5FFF7FFF9FFFBFFFDFFFF00010003",
		INIT_55=>X"FFFFFFFDFFFBFFFAFFF8FFF6FFF4FFF3FFF1FFF0FFEFFFEEFFEEFFEDFFEDFFED",
		INIT_56=>X"001100110011001100110010000F000E000D000C000A00090007000500030001",
		INIT_57=>X"FFFBFFFCFFFE000000020004000600070009000B000C000D000E000F00100011",
		INIT_58=>X"FFF0FFEFFFEFFFEFFFEEFFEEFFEFFFEFFFF0FFF1FFF2FFF3FFF4FFF6FFF7FFF9",
		INIT_59=>X"000900070005000400020000FFFEFFFDFFFBFFF9FFF7FFF6FFF4FFF3FFF2FFF1",
		INIT_5A=>X"000C000D000E000F000F00100010001000100010000F000E000E000D000B000A",
		INIT_5B=>X"FFF3FFF4FFF5FFF7FFF8FFFAFFFCFFFDFFFF000100030004000600080009000B",
		INIT_5C=>X"FFF7FFF6FFF4FFF3FFF2FFF1FFF0FFF0FFEFFFEFFFEFFFEFFFF0FFF0FFF1FFF2",
		INIT_5D=>X"000E000E000D000C000A000900080006000400030001FFFFFFFEFFFCFFFAFFF9",
		INIT_5E=>X"0004000500070008000A000B000C000D000E000F000F000F00100010000F000F",
		INIT_5F=>X"FFF0FFF0FFF0FFF1FFF2FFF3FFF4FFF5FFF6FFF8FFF9FFFBFFFDFFFE00000002",
		INIT_60=>X"0000FFFEFFFDFFFBFFF9FFF8FFF6FFF5FFF4FFF3FFF2FFF1FFF0FFF0FFF0FFF0",
		INIT_61=>X"000F00100010000F000F000F000E000D000C000B000A00080007000500040002",
		INIT_62=>X"FFFAFFFCFFFEFFFF000100030004000600080009000A000C000D000E000E000F",
		INIT_63=>X"FFF1FFF0FFF0FFEFFFEFFFEFFFEFFFF0FFF0FFF1FFF2FFF3FFF4FFF6FFF7FFF9",
		INIT_64=>X"000900080006000400030001FFFFFFFDFFFCFFFAFFF8FFF7FFF5FFF4FFF3FFF2",
		INIT_65=>X"000B000D000E000E000F00100010001000100010000F000F000E000D000C000B",
		INIT_66=>X"FFF2FFF3FFF4FFF6FFF7FFF9FFFBFFFDFFFE000000020004000500070009000A",
		INIT_67=>X"FFF7FFF6FFF4FFF3FFF2FFF1FFF0FFEFFFEFFFEEFFEEFFEFFFEFFFEFFFF0FFF1",
		INIT_68=>X"0010000F000E000D000C000B000900070006000400020000FFFEFFFCFFFBFFF9",
		INIT_69=>X"0003000500070009000A000C000D000E000F0010001100110011001100110011",
		INIT_6A=>X"FFEDFFEDFFEEFFEEFFEFFFF0FFF1FFF3FFF4FFF6FFF8FFFAFFFBFFFDFFFF0001",
		INIT_6B=>X"0001FFFFFFFDFFFBFFF9FFF7FFF5FFF4FFF2FFF1FFF0FFEFFFEEFFEDFFEDFFED",
		INIT_6C=>X"00130013001300130013001200120011000F000E000D000B0009000700050003",
		INIT_6D=>X"FFF8FFFAFFFCFFFE00000003000500070009000B000C000E000F001000110012",
		INIT_6E=>X"FFEDFFECFFEBFFEBFFEAFFEAFFEAFFEBFFECFFECFFEEFFEFFFF0FFF2FFF4FFF6",
		INIT_6F=>X"000E000C000A0007000500030000FFFEFFFCFFF9FFF7FFF5FFF3FFF1FFF0FFEE",
		INIT_70=>X"0010001100130014001500160016001700170016001600150014001300110010",
		INIT_71=>X"FFEBFFECFFEEFFF0FFF3FFF5FFF8FFFAFFFDFFFF0002000500070009000C000E",
		INIT_72=>X"FFF4FFF1FFEFFFEDFFEBFFEAFFE8FFE7FFE6FFE6FFE6FFE6FFE6FFE7FFE8FFE9",
		INIT_73=>X"001B001A00180016001400120010000D000A000800050002FFFFFFFCFFF9FFF6",
		INIT_74=>X"00040008000B000E00100013001500170019001A001B001C001C001D001C001C",
		INIT_75=>X"FFDEFFDEFFDFFFE0FFE2FFE3FFE6FFE8FFEBFFEDFFF1FFF4FFF7FFFAFFFE0001",
		INIT_76=>X"00050001FFFDFFF9FFF5FFF2FFEEFFEBFFE8FFE6FFE3FFE1FFE0FFDFFFDEFFDE",
		INIT_77=>X"002700280028002800270026002500230020001E001B001800140010000D0009",
		INIT_78=>X"FFECFFF1FFF5FFFAFFFF00040009000D001200160019001D0020002200240026",
		INIT_79=>X"FFD2FFCFFFCEFFCCFFCCFFCCFFCCFFCDFFCFFFD1FFD4FFD7FFDAFFDEFFE3FFE7",
		INIT_7A=>X"002B0025001F00180012000B0005FFFEFFF8FFF2FFECFFE6FFE1FFDDFFD8FFD5",
		INIT_7B=>X"00330039003D004100440046004800480048004600440042003E003A00350030",
		INIT_7C=>X"FFA4FFADFFB5FFBFFFC8FFD2FFDCFFE7FFF1FFFB0004000D0016001E0026002D",
		INIT_7D=>X"FFC2FFB5FFA9FF9FFF97FF91FF8BFF88FF86FF86FF86FF89FF8CFF91FF96FF9D",
		INIT_7E=>X"0129010F00F400DA00C000A6008D0074005C0044002E00190004FFF2FFE0FFD0",
		INIT_7F=>X"022E022B0226021E0215020A01FC01ED01DC01CA01B601A1018B0173015B0142",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_05,
		DOPADOP=>dopadop_05,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_06: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"00000FFFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF000000000000000",
		INITP_01=>X"00000000003FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFC000000000",
		INITP_02=>X"FC00000000000000FFFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF0000",
		INITP_03=>X"FFFFFFF000000000000003FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFF",
		INITP_04=>X"FFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFF000000000000003FFFFFFF",
		INITP_05=>X"0003FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFFC00000000000000FF",
		INITP_06=>X"000000000FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFF00000000000",
		INITP_07=>X"000000000000003FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFFC00000",
		INITP_08=>X"0003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000000",
		INITP_09=>X"00000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC000000",
		INITP_0A=>X"F0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF000",
		INITP_0B=>X"FFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF",
		INITP_0C=>X"FFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFF",
		INITP_0D=>X"003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003F",
		INITP_0E=>X"000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF00000000",
		INITP_0F=>X"0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000",
		INIT_00=>X"015B0173018B01A101B601CA01DC01ED01FC020A0215021E0226022B022E0230",
		INIT_01=>X"FFE0FFF200040019002E0044005C0074008D00A600C000DA00F4010F01290142",
		INIT_02=>X"FF96FF91FF8CFF89FF86FF86FF86FF88FF8BFF91FF97FF9FFFA9FFB5FFC2FFD0",
		INIT_03=>X"0026001E0016000D0004FFFBFFF1FFE7FFDCFFD2FFC8FFBFFFB5FFADFFA4FF9D",
		INIT_04=>X"0035003A003E004200440046004800480048004600440041003D00390033002D",
		INIT_05=>X"FFD8FFDDFFE1FFE6FFECFFF2FFF8FFFE0005000B00120018001F0025002B0030",
		INIT_06=>X"FFE3FFDEFFDAFFD7FFD4FFD1FFCFFFCDFFCCFFCCFFCCFFCCFFCEFFCFFFD2FFD5",
		INIT_07=>X"002400220020001D001900160012000D00090004FFFFFFFAFFF5FFF1FFECFFE7",
		INIT_08=>X"000D001000140018001B001E0020002300250026002700280028002800270026",
		INIT_09=>X"FFDEFFDFFFE0FFE1FFE3FFE6FFE8FFEBFFEEFFF2FFF5FFF9FFFD000100050009",
		INIT_0A=>X"FFFEFFFAFFF7FFF4FFF1FFEDFFEBFFE8FFE6FFE3FFE2FFE0FFDFFFDEFFDEFFDE",
		INIT_0B=>X"001C001D001C001C001B001A00190017001500130010000E000B000800040001",
		INIT_0C=>X"FFF9FFFCFFFF000200050008000A000D00100012001400160018001A001B001C",
		INIT_0D=>X"FFE8FFE7FFE6FFE6FFE6FFE6FFE6FFE7FFE8FFEAFFEBFFEDFFEFFFF1FFF4FFF6",
		INIT_0E=>X"000C0009000700050002FFFFFFFDFFFAFFF8FFF5FFF3FFF0FFEEFFECFFEBFFE9",
		INIT_0F=>X"001100130014001500160016001700170016001600150014001300110010000E",
		INIT_10=>X"FFF0FFF1FFF3FFF5FFF7FFF9FFFCFFFE0000000300050007000A000C000E0010",
		INIT_11=>X"FFF4FFF2FFF0FFEFFFEEFFECFFECFFEBFFEAFFEAFFEAFFEBFFEBFFECFFEDFFEE",
		INIT_12=>X"00110010000F000E000C000B00090007000500030000FFFEFFFCFFFAFFF8FFF6",
		INIT_13=>X"000500070009000B000D000E000F001100120012001300130013001300130012",
		INIT_14=>X"FFEDFFEDFFEEFFEFFFF0FFF1FFF2FFF4FFF5FFF7FFF9FFFBFFFDFFFF00010003",
		INIT_15=>X"FFFFFFFDFFFBFFFAFFF8FFF6FFF4FFF3FFF1FFF0FFEFFFEEFFEEFFEDFFEDFFED",
		INIT_16=>X"001100110011001100110010000F000E000D000C000A00090007000500030001",
		INIT_17=>X"FFFBFFFCFFFE000000020004000600070009000B000C000D000E000F00100011",
		INIT_18=>X"FFF0FFEFFFEFFFEFFFEEFFEEFFEFFFEFFFF0FFF1FFF2FFF3FFF4FFF6FFF7FFF9",
		INIT_19=>X"000900070005000400020000FFFEFFFDFFFBFFF9FFF7FFF6FFF4FFF3FFF2FFF1",
		INIT_1A=>X"000C000D000E000F000F00100010001000100010000F000E000E000D000B000A",
		INIT_1B=>X"FFF3FFF4FFF5FFF7FFF8FFFAFFFCFFFDFFFF000100030004000600080009000B",
		INIT_1C=>X"FFF7FFF6FFF4FFF3FFF2FFF1FFF0FFF0FFEFFFEFFFEFFFEFFFF0FFF0FFF1FFF2",
		INIT_1D=>X"000E000E000D000C000A000900080006000400030001FFFFFFFEFFFCFFFAFFF9",
		INIT_1E=>X"0004000500070008000A000B000C000D000E000F000F000F00100010000F000F",
		INIT_1F=>X"FFF0FFF0FFF0FFF1FFF2FFF3FFF4FFF5FFF6FFF8FFF9FFFBFFFDFFFE00000002",
		INIT_20=>X"0000FFFEFFFDFFFBFFF9FFF8FFF6FFF5FFF4FFF3FFF2FFF1FFF0FFF0FFF0FFF0",
		INIT_21=>X"000F00100010000F000F000F000E000D000C000B000A00080007000500040002",
		INIT_22=>X"FFFAFFFCFFFEFFFF000100030004000600080009000A000C000D000E000E000F",
		INIT_23=>X"FFF1FFF0FFF0FFEFFFEFFFEFFFEFFFF0FFF0FFF1FFF2FFF3FFF4FFF6FFF7FFF9",
		INIT_24=>X"000900080006000400030001FFFFFFFDFFFCFFFAFFF8FFF7FFF5FFF4FFF3FFF2",
		INIT_25=>X"000B000D000E000E000F00100010001000100010000F000F000E000D000C000B",
		INIT_26=>X"FFF2FFF3FFF4FFF6FFF7FFF9FFFBFFFDFFFE000000020004000500070009000A",
		INIT_27=>X"FFF7FFF6FFF4FFF3FFF2FFF1FFF0FFEFFFEFFFEEFFEEFFEFFFEFFFEFFFF0FFF1",
		INIT_28=>X"0010000F000E000D000C000B000900070006000400020000FFFEFFFCFFFBFFF9",
		INIT_29=>X"0003000500070009000A000C000D000E000F0010001100110011001100110011",
		INIT_2A=>X"FFEDFFEDFFEEFFEEFFEFFFF0FFF1FFF3FFF4FFF6FFF8FFFAFFFBFFFDFFFF0001",
		INIT_2B=>X"0001FFFFFFFDFFFBFFF9FFF7FFF5FFF4FFF2FFF1FFF0FFEFFFEEFFEDFFEDFFED",
		INIT_2C=>X"00130013001300130013001200120011000F000E000D000B0009000700050003",
		INIT_2D=>X"FFF8FFFAFFFCFFFE00000003000500070009000B000C000E000F001000110012",
		INIT_2E=>X"FFEDFFECFFEBFFEBFFEAFFEAFFEAFFEBFFECFFECFFEEFFEFFFF0FFF2FFF4FFF6",
		INIT_2F=>X"000E000C000A0007000500030000FFFEFFFCFFF9FFF7FFF5FFF3FFF1FFF0FFEE",
		INIT_30=>X"0010001100130014001500160016001700170016001600150014001300110010",
		INIT_31=>X"FFEBFFECFFEEFFF0FFF3FFF5FFF8FFFAFFFDFFFF0002000500070009000C000E",
		INIT_32=>X"FFF4FFF1FFEFFFEDFFEBFFEAFFE8FFE7FFE6FFE6FFE6FFE6FFE6FFE7FFE8FFE9",
		INIT_33=>X"001B001A00180016001400120010000D000A000800050002FFFFFFFCFFF9FFF6",
		INIT_34=>X"00040008000B000E00100013001500170019001A001B001C001C001D001C001C",
		INIT_35=>X"FFDEFFDEFFDFFFE0FFE2FFE3FFE6FFE8FFEBFFEDFFF1FFF4FFF7FFFAFFFE0001",
		INIT_36=>X"00050001FFFDFFF9FFF5FFF2FFEEFFEBFFE8FFE6FFE3FFE1FFE0FFDFFFDEFFDE",
		INIT_37=>X"002700280028002800270026002500230020001E001B001800140010000D0009",
		INIT_38=>X"FFECFFF1FFF5FFFAFFFF00040009000D001200160019001D0020002200240026",
		INIT_39=>X"FFD2FFCFFFCEFFCCFFCCFFCCFFCCFFCDFFCFFFD1FFD4FFD7FFDAFFDEFFE3FFE7",
		INIT_3A=>X"002B0025001F00180012000B0005FFFEFFF8FFF2FFECFFE6FFE1FFDDFFD8FFD5",
		INIT_3B=>X"00330039003D004100440046004800480048004600440042003E003A00350030",
		INIT_3C=>X"FFA4FFADFFB5FFBFFFC8FFD2FFDCFFE7FFF1FFFB0004000D0016001E0026002D",
		INIT_3D=>X"FFC2FFB5FFA9FF9FFF97FF91FF8BFF88FF86FF86FF86FF89FF8CFF91FF96FF9D",
		INIT_3E=>X"0129010F00F400DA00C000A6008D0074005C0044002E00190004FFF2FFE0FFD0",
		INIT_3F=>X"022E022B0226021E0215020A01FC01ED01DC01CA01B601A1018B0173015B0142",
		INIT_40=>X"00F8012F0166019E01D40209023B026B029602BD02DF02FB03120322032C0330",
		INIT_41=>X"FF59FF51FF4EFF4FFF55FF5FFF6EFF82FF9BFFB9FFDC0003002E005C008E00C2",
		INIT_42=>X"0061005A004F0043003400230010FFFCFFE7FFD2FFBDFFA8FF94FF81FF71FF63",
		INIT_43=>X"FFDDFFE8FFF500030011001E002C003900450050005900600065006800680066",
		INIT_44=>X"FFF2FFE8FFDEFFD4FFCCFFC4FFBEFFB9FFB6FFB4FFB5FFB7FFBBFFC1FFC9FFD2",
		INIT_45=>X"0029002F003400370039003A003A00370034002F00290022001900100006FFFC",
		INIT_46=>X"FFD0FFCFFFD0FFD2FFD5FFD9FFDEFFE4FFEBFFF3FFFB0003000B0013001B0022",
		INIT_47=>X"00230020001B00160010000A0003FFFCFFF5FFEEFFE8FFE2FFDDFFD8FFD4FFD1",
		INIT_48=>X"FFF1FFF7FFFD00030009000F00140019001E0022002500270028002900280026",
		INIT_49=>X"FFF7FFF2FFEDFFE8FFE5FFE1FFDFFFDDFFDCFFDCFFDCFFDEFFE0FFE4FFE8FFEC",
		INIT_4A=>X"0018001B001D001F001F001F001F001D001B001800140010000C00070001FFFC",
		INIT_4B=>X"FFE3FFE3FFE3FFE5FFE7FFEAFFEDFFF1FFF5FFF9FFFE00030008000C00100014",
		INIT_4C=>X"001600130010000D000900050000FFFCFFF8FFF4FFF0FFECFFE9FFE7FFE5FFE3",
		INIT_4D=>X"FFF7FFFBFFFF00030007000B000E00110014001700180019001A001A00190018",
		INIT_4E=>X"FFF8FFF5FFF2FFEFFFECFFEAFFE8FFE7FFE7FFE7FFE8FFE9FFEBFFEDFFF0FFF4",
		INIT_4F=>X"0012001400150016001600160016001400120010000D000A000700030000FFFC",
		INIT_50=>X"FFEAFFEAFFEBFFECFFEEFFF0FFF3FFF6FFF9FFFC000000030006000A000D0010",
		INIT_51=>X"0010000E000B000900060002FFFFFFFCFFF9FFF6FFF3FFF0FFEEFFECFFEBFFEA",
		INIT_52=>X"FFFAFFFD0000000300060009000C000E00100012001300140014001400130012",
		INIT_53=>X"FFF9FFF6FFF4FFF1FFEFFFEEFFEDFFECFFECFFECFFEDFFEEFFF0FFF2FFF4FFF7",
		INIT_54=>X"000F0011001200120012001200110010000E000C000A000700050002FFFFFFFC",
		INIT_55=>X"FFEDFFEEFFEFFFF0FFF1FFF3FFF6FFF8FFFBFFFE0000000300060009000B000D",
		INIT_56=>X"000D000B0009000700040001FFFEFFFCFFF9FFF6FFF4FFF2FFF0FFEFFFEEFFED",
		INIT_57=>X"FFFBFFFE0001000400060009000B000D000E001000110011001100110010000F",
		INIT_58=>X"FFF9FFF6FFF4FFF2FFF1FFF0FFEFFFEEFFEEFFEFFFF0FFF1FFF2FFF4FFF6FFF9",
		INIT_59=>X"000E000F0010001000100010000F000E000C000A0008000600030001FFFEFFFB",
		INIT_5A=>X"FFEFFFF0FFF0FFF2FFF3FFF5FFF7FFFAFFFCFFFF0001000400060009000B000C",
		INIT_5B=>X"000B000A0008000500030000FFFEFFFBFFF9FFF6FFF4FFF3FFF1FFF0FFEFFFEF",
		INIT_5C=>X"FFFCFFFF0002000400060009000B000C000E000F000F00100010000F000E000D",
		INIT_5D=>X"FFF8FFF6FFF4FFF3FFF1FFF0FFF0FFEFFFF0FFF0FFF1FFF2FFF4FFF6FFF8FFFA",
		INIT_5E=>X"000E000F000F0010000F000F000E000D000B00090007000500020000FFFDFFFB",
		INIT_5F=>X"FFF0FFF0FFF1FFF3FFF4FFF6FFF8FFFAFFFDFFFF0002000400070009000B000C",
		INIT_60=>X"000B0009000700040002FFFFFFFDFFFAFFF8FFF6FFF4FFF3FFF1FFF0FFF0FFF0",
		INIT_61=>X"FFFD00000002000500070009000B000D000E000F000F0010000F000F000E000C",
		INIT_62=>X"FFF8FFF6FFF4FFF2FFF1FFF0FFF0FFEFFFF0FFF0FFF1FFF3FFF4FFF6FFF8FFFB",
		INIT_63=>X"000E000F00100010000F000F000E000C000B0009000600040002FFFFFFFCFFFA",
		INIT_64=>X"FFEFFFF0FFF1FFF3FFF4FFF6FFF9FFFBFFFE0000000300050008000A000B000D",
		INIT_65=>X"000B0009000600040001FFFFFFFCFFFAFFF7FFF5FFF3FFF2FFF0FFF0FFEFFFEF",
		INIT_66=>X"FFFE0001000300060008000A000C000E000F0010001000100010000F000E000C",
		INIT_67=>X"FFF6FFF4FFF2FFF1FFF0FFEFFFEEFFEEFFEFFFF0FFF1FFF2FFF4FFF6FFF9FFFB",
		INIT_68=>X"001000110011001100110010000E000D000B0009000600040001FFFEFFFBFFF9",
		INIT_69=>X"FFEEFFEFFFF0FFF2FFF4FFF6FFF9FFFCFFFE0001000400070009000B000D000F",
		INIT_6A=>X"000B0009000600030000FFFEFFFBFFF8FFF6FFF3FFF1FFF0FFEFFFEEFFEDFFED",
		INIT_6B=>X"FFFF000200050007000A000C000E0010001100120012001200120011000F000D",
		INIT_6C=>X"FFF4FFF2FFF0FFEEFFEDFFECFFECFFECFFEDFFEEFFEFFFF1FFF4FFF6FFF9FFFC",
		INIT_6D=>X"0013001400140014001300120010000E000C0009000600030000FFFDFFFAFFF7",
		INIT_6E=>X"FFEBFFECFFEEFFF0FFF3FFF6FFF9FFFCFFFF000200060009000B000E00100012",
		INIT_6F=>X"000D000A000600030000FFFCFFF9FFF6FFF3FFF0FFEEFFECFFEBFFEAFFEAFFEA",
		INIT_70=>X"000000030007000A000D00100012001400160016001600160015001400120010",
		INIT_71=>X"FFF0FFEDFFEBFFE9FFE8FFE7FFE7FFE7FFE8FFEAFFECFFEFFFF2FFF5FFF8FFFC",
		INIT_72=>X"0019001A001A00190018001700140011000E000B00070003FFFFFFFBFFF7FFF4",
		INIT_73=>X"FFE5FFE7FFE9FFECFFF0FFF4FFF8FFFC000000050009000D0010001300160018",
		INIT_74=>X"0010000C00080003FFFEFFF9FFF5FFF1FFEDFFEAFFE7FFE5FFE3FFE3FFE3FFE3",
		INIT_75=>X"00010007000C001000140018001B001D001F001F001F001F001D001B00180014",
		INIT_76=>X"FFE8FFE4FFE0FFDEFFDCFFDCFFDCFFDDFFDFFFE1FFE5FFE8FFEDFFF2FFF7FFFC",
		INIT_77=>X"002800290028002700250022001E00190014000F00090003FFFDFFF7FFF1FFEC",
		INIT_78=>X"FFD4FFD8FFDDFFE2FFE8FFEEFFF5FFFC0003000A00100016001B002000230026",
		INIT_79=>X"001B0013000B0003FFFBFFF3FFEBFFE4FFDEFFD9FFD5FFD2FFD0FFCFFFD0FFD1",
		INIT_7A=>X"00060010001900220029002F00340037003A003A003900370034002F00290022",
		INIT_7B=>X"FFC9FFC1FFBBFFB7FFB5FFB4FFB6FFB9FFBEFFC4FFCCFFD4FFDEFFE8FFF2FFFC",
		INIT_7C=>X"00680068006500600059005000450039002C001E00110003FFF5FFE8FFDDFFD2",
		INIT_7D=>X"FF71FF81FF94FFA8FFBDFFD2FFE7FFFC0010002300340043004F005A00610066",
		INIT_7E=>X"008E005C002E0003FFDCFFB9FF9BFF82FF6EFF5FFF55FF4FFF4EFF51FF59FF63",
		INIT_7F=>X"032C0322031202FB02DF02BD0296026B023B020901D4019E0166012F00F800C2",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_06,
		DOPADOP=>dopadop_06,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_07: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"0003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000000",
		INITP_01=>X"00000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC000000",
		INITP_02=>X"F0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF000",
		INITP_03=>X"FFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF",
		INITP_04=>X"FFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFF",
		INITP_05=>X"003FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000003F",
		INITP_06=>X"000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF00000000",
		INITP_07=>X"0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000",
		INITP_08=>X"000000FFFFFFFC0000003FFFFFFC0000000FFFFFFF00000003FFFFFFC0000000",
		INITP_09=>X"FFFFF00000003FFFFFFC0000000FFFFFFF0000000FFFFFFFC0000003FFFFFFF0",
		INITP_0A=>X"00003FFFFFFC0000003FFFFFFF0000000FFFFFFFC0000003FFFFFFC0000000FF",
		INITP_0B=>X"FFFC0000003FFFFFFF0000000FFFFFFF00000003FFFFFFC0000000FFFFFFF000",
		INITP_0C=>X"003FFFFFFC0000000FFFFFFF00000003FFFFFFC0000003FFFFFFF0000000FFFF",
		INITP_0D=>X"FC0000000FFFFFFF0000000FFFFFFFC0000003FFFFFFF0000000FFFFFFF00000",
		INITP_0E=>X"3FFFFFFF0000000FFFFFFFC0000003FFFFFFC0000000FFFFFFF00000003FFFFF",
		INITP_0F=>X"0000000FFFFFFF00000003FFFFFFC0000000FFFFFFF0000000FFFFFFFC000000",
		INIT_00=>X"00F8012F0166019E01D40209023B026B029602BD02DF02FB03120322032C0330",
		INIT_01=>X"FF59FF51FF4EFF4FFF55FF5FFF6EFF82FF9BFFB9FFDC0003002E005C008E00C2",
		INIT_02=>X"0061005A004F0043003400230010FFFCFFE7FFD2FFBDFFA8FF94FF81FF71FF63",
		INIT_03=>X"FFDDFFE8FFF500030011001E002C003900450050005900600065006800680066",
		INIT_04=>X"FFF2FFE8FFDEFFD4FFCCFFC4FFBEFFB9FFB6FFB4FFB5FFB7FFBBFFC1FFC9FFD2",
		INIT_05=>X"0029002F003400370039003A003A00370034002F00290022001900100006FFFC",
		INIT_06=>X"FFD0FFCFFFD0FFD2FFD5FFD9FFDEFFE4FFEBFFF3FFFB0003000B0013001B0022",
		INIT_07=>X"00230020001B00160010000A0003FFFCFFF5FFEEFFE8FFE2FFDDFFD8FFD4FFD1",
		INIT_08=>X"FFF1FFF7FFFD00030009000F00140019001E0022002500270028002900280026",
		INIT_09=>X"FFF7FFF2FFEDFFE8FFE5FFE1FFDFFFDDFFDCFFDCFFDCFFDEFFE0FFE4FFE8FFEC",
		INIT_0A=>X"0018001B001D001F001F001F001F001D001B001800140010000C00070001FFFC",
		INIT_0B=>X"FFE3FFE3FFE3FFE5FFE7FFEAFFEDFFF1FFF5FFF9FFFE00030008000C00100014",
		INIT_0C=>X"001600130010000D000900050000FFFCFFF8FFF4FFF0FFECFFE9FFE7FFE5FFE3",
		INIT_0D=>X"FFF7FFFBFFFF00030007000B000E00110014001700180019001A001A00190018",
		INIT_0E=>X"FFF8FFF5FFF2FFEFFFECFFEAFFE8FFE7FFE7FFE7FFE8FFE9FFEBFFEDFFF0FFF4",
		INIT_0F=>X"0012001400150016001600160016001400120010000D000A000700030000FFFC",
		INIT_10=>X"FFEAFFEAFFEBFFECFFEEFFF0FFF3FFF6FFF9FFFC000000030006000A000D0010",
		INIT_11=>X"0010000E000B000900060002FFFFFFFCFFF9FFF6FFF3FFF0FFEEFFECFFEBFFEA",
		INIT_12=>X"FFFAFFFD0000000300060009000C000E00100012001300140014001400130012",
		INIT_13=>X"FFF9FFF6FFF4FFF1FFEFFFEEFFEDFFECFFECFFECFFEDFFEEFFF0FFF2FFF4FFF7",
		INIT_14=>X"000F0011001200120012001200110010000E000C000A000700050002FFFFFFFC",
		INIT_15=>X"FFEDFFEEFFEFFFF0FFF1FFF3FFF6FFF8FFFBFFFE0000000300060009000B000D",
		INIT_16=>X"000D000B0009000700040001FFFEFFFCFFF9FFF6FFF4FFF2FFF0FFEFFFEEFFED",
		INIT_17=>X"FFFBFFFE0001000400060009000B000D000E001000110011001100110010000F",
		INIT_18=>X"FFF9FFF6FFF4FFF2FFF1FFF0FFEFFFEEFFEEFFEFFFF0FFF1FFF2FFF4FFF6FFF9",
		INIT_19=>X"000E000F0010001000100010000F000E000C000A0008000600030001FFFEFFFB",
		INIT_1A=>X"FFEFFFF0FFF0FFF2FFF3FFF5FFF7FFFAFFFCFFFF0001000400060009000B000C",
		INIT_1B=>X"000B000A0008000500030000FFFEFFFBFFF9FFF6FFF4FFF3FFF1FFF0FFEFFFEF",
		INIT_1C=>X"FFFCFFFF0002000400060009000B000C000E000F000F00100010000F000E000D",
		INIT_1D=>X"FFF8FFF6FFF4FFF3FFF1FFF0FFF0FFEFFFF0FFF0FFF1FFF2FFF4FFF6FFF8FFFA",
		INIT_1E=>X"000E000F000F0010000F000F000E000D000B00090007000500020000FFFDFFFB",
		INIT_1F=>X"FFF0FFF0FFF1FFF3FFF4FFF6FFF8FFFAFFFDFFFF0002000400070009000B000C",
		INIT_20=>X"000B0009000700040002FFFFFFFDFFFAFFF8FFF6FFF4FFF3FFF1FFF0FFF0FFF0",
		INIT_21=>X"FFFD00000002000500070009000B000D000E000F000F0010000F000F000E000C",
		INIT_22=>X"FFF8FFF6FFF4FFF2FFF1FFF0FFF0FFEFFFF0FFF0FFF1FFF3FFF4FFF6FFF8FFFB",
		INIT_23=>X"000E000F00100010000F000F000E000C000B0009000600040002FFFFFFFCFFFA",
		INIT_24=>X"FFEFFFF0FFF1FFF3FFF4FFF6FFF9FFFBFFFE0000000300050008000A000B000D",
		INIT_25=>X"000B0009000600040001FFFFFFFCFFFAFFF7FFF5FFF3FFF2FFF0FFF0FFEFFFEF",
		INIT_26=>X"FFFE0001000300060008000A000C000E000F0010001000100010000F000E000C",
		INIT_27=>X"FFF6FFF4FFF2FFF1FFF0FFEFFFEEFFEEFFEFFFF0FFF1FFF2FFF4FFF6FFF9FFFB",
		INIT_28=>X"001000110011001100110010000E000D000B0009000600040001FFFEFFFBFFF9",
		INIT_29=>X"FFEEFFEFFFF0FFF2FFF4FFF6FFF9FFFCFFFE0001000400070009000B000D000F",
		INIT_2A=>X"000B0009000600030000FFFEFFFBFFF8FFF6FFF3FFF1FFF0FFEFFFEEFFEDFFED",
		INIT_2B=>X"FFFF000200050007000A000C000E0010001100120012001200120011000F000D",
		INIT_2C=>X"FFF4FFF2FFF0FFEEFFEDFFECFFECFFECFFEDFFEEFFEFFFF1FFF4FFF6FFF9FFFC",
		INIT_2D=>X"0013001400140014001300120010000E000C0009000600030000FFFDFFFAFFF7",
		INIT_2E=>X"FFEBFFECFFEEFFF0FFF3FFF6FFF9FFFCFFFF000200060009000B000E00100012",
		INIT_2F=>X"000D000A000600030000FFFCFFF9FFF6FFF3FFF0FFEEFFECFFEBFFEAFFEAFFEA",
		INIT_30=>X"000000030007000A000D00100012001400160016001600160015001400120010",
		INIT_31=>X"FFF0FFEDFFEBFFE9FFE8FFE7FFE7FFE7FFE8FFEAFFECFFEFFFF2FFF5FFF8FFFC",
		INIT_32=>X"0019001A001A00190018001700140011000E000B00070003FFFFFFFBFFF7FFF4",
		INIT_33=>X"FFE5FFE7FFE9FFECFFF0FFF4FFF8FFFC000000050009000D0010001300160018",
		INIT_34=>X"0010000C00080003FFFEFFF9FFF5FFF1FFEDFFEAFFE7FFE5FFE3FFE3FFE3FFE3",
		INIT_35=>X"00010007000C001000140018001B001D001F001F001F001F001D001B00180014",
		INIT_36=>X"FFE8FFE4FFE0FFDEFFDCFFDCFFDCFFDDFFDFFFE1FFE5FFE8FFEDFFF2FFF7FFFC",
		INIT_37=>X"002800290028002700250022001E00190014000F00090003FFFDFFF7FFF1FFEC",
		INIT_38=>X"FFD4FFD8FFDDFFE2FFE8FFEEFFF5FFFC0003000A00100016001B002000230026",
		INIT_39=>X"001B0013000B0003FFFBFFF3FFEBFFE4FFDEFFD9FFD5FFD2FFD0FFCFFFD0FFD1",
		INIT_3A=>X"00060010001900220029002F00340037003A003A003900370034002F00290022",
		INIT_3B=>X"FFC9FFC1FFBBFFB7FFB5FFB4FFB6FFB9FFBEFFC4FFCCFFD4FFDEFFE8FFF2FFFC",
		INIT_3C=>X"00680068006500600059005000450039002C001E00110003FFF5FFE8FFDDFFD2",
		INIT_3D=>X"FF71FF81FF94FFA8FFBDFFD2FFE7FFFC0010002300340043004F005A00610066",
		INIT_3E=>X"008E005C002E0003FFDCFFB9FF9BFF82FF6EFF5FFF55FF4FFF4EFF51FF59FF63",
		INIT_3F=>X"032C0322031202FB02DF02BD0296026B023B020901D4019E0166012F00F800C2",
		INIT_40=>X"FFD40022007A00DA014101AC0218028202E80347039C03E50420044C04670470",
		INIT_41=>X"004C002B0006FFDDFFB4FF8BFF64FF42FF27FF13FF09FF0BFF19FF34FF5CFF92",
		INIT_42=>X"FFAFFFC0FFD5FFED00070021003C0055006B007D008A00910091008A007C0067",
		INIT_43=>X"004C00440038002A00190006FFF2FFDEFFCBFFBAFFABFFA0FF99FF97FF9AFFA2",
		INIT_44=>X"FFBDFFBFFFC4FFCCFFD6FFE3FFF2000100110021002F003C0046004D00500050",
		INIT_45=>X"0035003800380035002F0028001E00120006FFF8FFEBFFDFFFD3FFCAFFC3FFBE",
		INIT_46=>X"FFD8FFD3FFD0FFCEFFCFFFD3FFD9FFE0FFE9FFF4FFFF000A0016002000290030",
		INIT_47=>X"0018001F00250029002B002B00290025001F0018000F0006FFFCFFF2FFE8FFE0",
		INIT_48=>X"FFF6FFEEFFE7FFE1FFDCFFD9FFD8FFD9FFDCFFE0FFE6FFEDFFF5FFFE00070010",
		INIT_49=>X"FFFD0004000C00120018001D0021002300230022001F001A0014000D0006FFFE",
		INIT_4A=>X"000C0006FFFFFFF8FFF2FFECFFE6FFE3FFE0FFDFFFDFFFE1FFE4FFE9FFEFFFF6",
		INIT_4B=>X"FFEBFFF0FFF6FFFC00030009000F00140018001C001D001E001D001B00170012",
		INIT_4C=>X"001800150010000B00060000FFFAFFF4FFEFFFEAFFE7FFE4FFE3FFE3FFE5FFE8",
		INIT_4D=>X"FFE6FFE8FFEAFFEDFFF1FFF6FFFC00010007000C001100150018001A001A001A",
		INIT_4E=>X"00170017001700150013000F000B00060001FFFBFFF6FFF1FFEDFFEAFFE8FFE6",
		INIT_4F=>X"FFECFFEAFFE9FFE9FFEAFFECFFEEFFF2FFF7FFFB00000005000A000F00120015",
		INIT_50=>X"000D0010001300150015001500140012000E000B00060001FFFDFFF8FFF3FFF0",
		INIT_51=>X"FFF9FFF5FFF1FFEEFFECFFEBFFEAFFEBFFEDFFEFFFF3FFF7FFFB000000040009",
		INIT_52=>X"FFFF00030007000B000F001100130014001400130011000E000A00060002FFFD",
		INIT_53=>X"00060002FFFEFFFAFFF6FFF3FFF0FFEEFFECFFECFFECFFEEFFF0FFF3FFF7FFFB",
		INIT_54=>X"FFF3FFF7FFFAFFFE00020006000A000D001000120012001200120010000D000A",
		INIT_55=>X"000F000D000A00070003FFFFFFFBFFF7FFF4FFF1FFEFFFEDFFEDFFEDFFEFFFF1",
		INIT_56=>X"FFEEFFEFFFF1FFF3FFF6FFFAFFFE000200050009000C000F0010001100120011",
		INIT_57=>X"001100110010000F000D000A000700030000FFFCFFF8FFF5FFF2FFF0FFEEFFEE",
		INIT_58=>X"FFF1FFEFFFEFFFEFFFEFFFF1FFF3FFF6FFFAFFFD000100050008000B000E0010",
		INIT_59=>X"000A000D000F001000100010000F000D000A000700040000FFFCFFF9FFF6FFF3",
		INIT_5A=>X"FFFAFFF6FFF4FFF1FFF0FFEFFFEFFFF0FFF1FFF3FFF6FFF9FFFD000000040007",
		INIT_5B=>X"000000030007000A000C000E000F00100010000F000D000A000700040001FFFD",
		INIT_5C=>X"00050001FFFEFFFAFFF7FFF4FFF2FFF0FFEFFFEFFFF0FFF1FFF3FFF6FFF9FFFC",
		INIT_5D=>X"FFF6FFF9FFFCFFFF000300060009000C000E000F0010000F000F000D000B0008",
		INIT_5E=>X"000D000B000800050002FFFEFFFBFFF8FFF5FFF2FFF1FFF0FFEFFFF0FFF1FFF3",
		INIT_5F=>X"FFF0FFF1FFF3FFF5FFF8FFFBFFFF000200060009000B000D000F000F000F000F",
		INIT_60=>X"000F000F000F000D000B000900060002FFFFFFFBFFF8FFF5FFF3FFF1FFF0FFF0",
		INIT_61=>X"FFF1FFF0FFEFFFF0FFF1FFF2FFF5FFF8FFFBFFFE000200050008000B000D000F",
		INIT_62=>X"000B000D000F000F0010000F000E000C000900060003FFFFFFFCFFF9FFF6FFF3",
		INIT_63=>X"FFF9FFF6FFF3FFF1FFF0FFEFFFEFFFF0FFF2FFF4FFF7FFFAFFFE000100050008",
		INIT_64=>X"000100040007000A000D000F00100010000F000E000C000A000700030000FFFC",
		INIT_65=>X"00040000FFFDFFF9FFF6FFF3FFF1FFF0FFEFFFEFFFF0FFF1FFF4FFF6FFFAFFFD",
		INIT_66=>X"FFF6FFF9FFFC000000040007000A000D000F001000100010000F000D000A0007",
		INIT_67=>X"000E000B000800050001FFFDFFFAFFF6FFF3FFF1FFEFFFEFFFEFFFEFFFF1FFF3",
		INIT_68=>X"FFEEFFF0FFF2FFF5FFF8FFFC000000030007000A000D000F0010001100110010",
		INIT_69=>X"001200110010000F000C000900050002FFFEFFFAFFF6FFF3FFF1FFEFFFEEFFEE",
		INIT_6A=>X"FFEFFFEDFFEDFFEDFFEFFFF1FFF4FFF7FFFBFFFF00030007000A000D000F0011",
		INIT_6B=>X"000D001000120012001200120010000D000A00060002FFFEFFFAFFF7FFF3FFF1",
		INIT_6C=>X"FFF7FFF3FFF0FFEEFFECFFECFFECFFEEFFF0FFF3FFF6FFFAFFFE00020006000A",
		INIT_6D=>X"00020006000A000E001100130014001400130011000F000B00070003FFFFFFFB",
		INIT_6E=>X"00040000FFFBFFF7FFF3FFEFFFEDFFEBFFEAFFEBFFECFFEEFFF1FFF5FFF9FFFD",
		INIT_6F=>X"FFF3FFF8FFFD00010006000B000E0012001400150015001500130010000D0009",
		INIT_70=>X"0012000F000A00050000FFFBFFF7FFF2FFEEFFECFFEAFFE9FFE9FFEAFFECFFF0",
		INIT_71=>X"FFE8FFEAFFEDFFF1FFF6FFFB00010006000B000F001300150017001700170015",
		INIT_72=>X"001A001A001800150011000C00070001FFFCFFF6FFF1FFEDFFEAFFE8FFE6FFE6",
		INIT_73=>X"FFE5FFE3FFE3FFE4FFE7FFEAFFEFFFF4FFFA00000006000B001000150018001A",
		INIT_74=>X"0017001B001D001E001D001C00180014000F00090003FFFCFFF6FFF0FFEBFFE8",
		INIT_75=>X"FFEFFFE9FFE4FFE1FFDFFFDFFFE0FFE3FFE6FFECFFF2FFF8FFFF0006000C0012",
		INIT_76=>X"0006000D0014001A001F0022002300230021001D00180012000C0004FFFDFFF6",
		INIT_77=>X"0007FFFEFFF5FFEDFFE6FFE0FFDCFFD9FFD8FFD9FFDCFFE1FFE7FFEEFFF6FFFE",
		INIT_78=>X"FFE8FFF2FFFC0006000F0018001F00250029002B002B00290025001F00180010",
		INIT_79=>X"002900200016000AFFFFFFF4FFE9FFE0FFD9FFD3FFCFFFCEFFD0FFD3FFD8FFE0",
		INIT_7A=>X"FFC3FFCAFFD3FFDFFFEBFFF800060012001E0028002F00350038003800350030",
		INIT_7B=>X"0050004D0046003C002F002100110001FFF2FFE3FFD6FFCCFFC4FFBFFFBDFFBE",
		INIT_7C=>X"FF9AFF97FF99FFA0FFABFFBAFFCBFFDEFFF200060019002A00380044004C0050",
		INIT_7D=>X"007C008A00910091008A007D006B0055003C00210007FFEDFFD5FFC0FFAFFFA2",
		INIT_7E=>X"FF5CFF34FF19FF0BFF09FF13FF27FF42FF64FF8BFFB4FFDD0006002B004C0067",
		INIT_7F=>X"0467044C042003E5039C034702E80282021801AC014100DA007A0022FFD4FF92",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_07,
		DOPADOP=>dopadop_07,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_08: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"000000FFFFFFFC0000003FFFFFFC0000000FFFFFFF00000003FFFFFFC0000000",
		INITP_01=>X"FFFFF00000003FFFFFFC0000000FFFFFFF0000000FFFFFFFC0000003FFFFFFF0",
		INITP_02=>X"00003FFFFFFC0000003FFFFFFF0000000FFFFFFFC0000003FFFFFFC0000000FF",
		INITP_03=>X"FFFC0000003FFFFFFF0000000FFFFFFF00000003FFFFFFC0000000FFFFFFF000",
		INITP_04=>X"003FFFFFFC0000000FFFFFFF00000003FFFFFFC0000003FFFFFFF0000000FFFF",
		INITP_05=>X"FC0000000FFFFFFF0000000FFFFFFFC0000003FFFFFFF0000000FFFFFFF00000",
		INITP_06=>X"3FFFFFFF0000000FFFFFFFC0000003FFFFFFC0000000FFFFFFF00000003FFFFF",
		INITP_07=>X"0000000FFFFFFF00000003FFFFFFC0000000FFFFFFF0000000FFFFFFFC000000",
		INITP_08=>X"000FFFFF00000FFFFF00000FFFFFC00003FFFFC00003FFFFC00003FFFFC00000",
		INITP_09=>X"F00000FFFFF00000FFFFFC00003FFFFC00003FFFFC00003FFFFC00000FFFFF00",
		INITP_0A=>X"FFFF000003FFFFC00003FFFFC00003FFFFC00003FFFFC00000FFFFF00000FFFF",
		INITP_0B=>X"003FFFFC00003FFFFC00003FFFFC00003FFFFF00000FFFFF00000FFFFF00000F",
		INITP_0C=>X"C00003FFFFC00003FFFFC00003FFFFF00000FFFFF00000FFFFF00000FFFFF000",
		INITP_0D=>X"FFFC00003FFFFC00000FFFFF00000FFFFF00000FFFFF00000FFFFF000003FFFF",
		INITP_0E=>X"03FFFFC00000FFFFF00000FFFFF00000FFFFF00000FFFFFC00003FFFFC00003F",
		INITP_0F=>X"00000FFFFF00000FFFFF00000FFFFF00000FFFFFC00003FFFFC00003FFFFC000",
		INIT_00=>X"FFD40022007A00DA014101AC0218028202E80347039C03E50420044C04670470",
		INIT_01=>X"004C002B0006FFDDFFB4FF8BFF64FF42FF27FF13FF09FF0BFF19FF34FF5CFF92",
		INIT_02=>X"FFAFFFC0FFD5FFED00070021003C0055006B007D008A00910091008A007C0067",
		INIT_03=>X"004C00440038002A00190006FFF2FFDEFFCBFFBAFFABFFA0FF99FF97FF9AFFA2",
		INIT_04=>X"FFBDFFBFFFC4FFCCFFD6FFE3FFF2000100110021002F003C0046004D00500050",
		INIT_05=>X"0035003800380035002F0028001E00120006FFF8FFEBFFDFFFD3FFCAFFC3FFBE",
		INIT_06=>X"FFD8FFD3FFD0FFCEFFCFFFD3FFD9FFE0FFE9FFF4FFFF000A0016002000290030",
		INIT_07=>X"0018001F00250029002B002B00290025001F0018000F0006FFFCFFF2FFE8FFE0",
		INIT_08=>X"FFF6FFEEFFE7FFE1FFDCFFD9FFD8FFD9FFDCFFE0FFE6FFEDFFF5FFFE00070010",
		INIT_09=>X"FFFD0004000C00120018001D0021002300230022001F001A0014000D0006FFFE",
		INIT_0A=>X"000C0006FFFFFFF8FFF2FFECFFE6FFE3FFE0FFDFFFDFFFE1FFE4FFE9FFEFFFF6",
		INIT_0B=>X"FFEBFFF0FFF6FFFC00030009000F00140018001C001D001E001D001B00170012",
		INIT_0C=>X"001800150010000B00060000FFFAFFF4FFEFFFEAFFE7FFE4FFE3FFE3FFE5FFE8",
		INIT_0D=>X"FFE6FFE8FFEAFFEDFFF1FFF6FFFC00010007000C001100150018001A001A001A",
		INIT_0E=>X"00170017001700150013000F000B00060001FFFBFFF6FFF1FFEDFFEAFFE8FFE6",
		INIT_0F=>X"FFECFFEAFFE9FFE9FFEAFFECFFEEFFF2FFF7FFFB00000005000A000F00120015",
		INIT_10=>X"000D0010001300150015001500140012000E000B00060001FFFDFFF8FFF3FFF0",
		INIT_11=>X"FFF9FFF5FFF1FFEEFFECFFEBFFEAFFEBFFEDFFEFFFF3FFF7FFFB000000040009",
		INIT_12=>X"FFFF00030007000B000F001100130014001400130011000E000A00060002FFFD",
		INIT_13=>X"00060002FFFEFFFAFFF6FFF3FFF0FFEEFFECFFECFFECFFEEFFF0FFF3FFF7FFFB",
		INIT_14=>X"FFF3FFF7FFFAFFFE00020006000A000D001000120012001200120010000D000A",
		INIT_15=>X"000F000D000A00070003FFFFFFFBFFF7FFF4FFF1FFEFFFEDFFEDFFEDFFEFFFF1",
		INIT_16=>X"FFEEFFEFFFF1FFF3FFF6FFFAFFFE000200050009000C000F0010001100120011",
		INIT_17=>X"001100110010000F000D000A000700030000FFFCFFF8FFF5FFF2FFF0FFEEFFEE",
		INIT_18=>X"FFF1FFEFFFEFFFEFFFEFFFF1FFF3FFF6FFFAFFFD000100050008000B000E0010",
		INIT_19=>X"000A000D000F001000100010000F000D000A000700040000FFFCFFF9FFF6FFF3",
		INIT_1A=>X"FFFAFFF6FFF4FFF1FFF0FFEFFFEFFFF0FFF1FFF3FFF6FFF9FFFD000000040007",
		INIT_1B=>X"000000030007000A000C000E000F00100010000F000D000A000700040001FFFD",
		INIT_1C=>X"00050001FFFEFFFAFFF7FFF4FFF2FFF0FFEFFFEFFFF0FFF1FFF3FFF6FFF9FFFC",
		INIT_1D=>X"FFF6FFF9FFFCFFFF000300060009000C000E000F0010000F000F000D000B0008",
		INIT_1E=>X"000D000B000800050002FFFEFFFBFFF8FFF5FFF2FFF1FFF0FFEFFFF0FFF1FFF3",
		INIT_1F=>X"FFF0FFF1FFF3FFF5FFF8FFFBFFFF000200060009000B000D000F000F000F000F",
		INIT_20=>X"000F000F000F000D000B000900060002FFFFFFFBFFF8FFF5FFF3FFF1FFF0FFF0",
		INIT_21=>X"FFF1FFF0FFEFFFF0FFF1FFF2FFF5FFF8FFFBFFFE000200050008000B000D000F",
		INIT_22=>X"000B000D000F000F0010000F000E000C000900060003FFFFFFFCFFF9FFF6FFF3",
		INIT_23=>X"FFF9FFF6FFF3FFF1FFF0FFEFFFEFFFF0FFF2FFF4FFF7FFFAFFFE000100050008",
		INIT_24=>X"000100040007000A000D000F00100010000F000E000C000A000700030000FFFC",
		INIT_25=>X"00040000FFFDFFF9FFF6FFF3FFF1FFF0FFEFFFEFFFF0FFF1FFF4FFF6FFFAFFFD",
		INIT_26=>X"FFF6FFF9FFFC000000040007000A000D000F001000100010000F000D000A0007",
		INIT_27=>X"000E000B000800050001FFFDFFFAFFF6FFF3FFF1FFEFFFEFFFEFFFEFFFF1FFF3",
		INIT_28=>X"FFEEFFF0FFF2FFF5FFF8FFFC000000030007000A000D000F0010001100110010",
		INIT_29=>X"001200110010000F000C000900050002FFFEFFFAFFF6FFF3FFF1FFEFFFEEFFEE",
		INIT_2A=>X"FFEFFFEDFFEDFFEDFFEFFFF1FFF4FFF7FFFBFFFF00030007000A000D000F0011",
		INIT_2B=>X"000D001000120012001200120010000D000A00060002FFFEFFFAFFF7FFF3FFF1",
		INIT_2C=>X"FFF7FFF3FFF0FFEEFFECFFECFFECFFEEFFF0FFF3FFF6FFFAFFFE00020006000A",
		INIT_2D=>X"00020006000A000E001100130014001400130011000F000B00070003FFFFFFFB",
		INIT_2E=>X"00040000FFFBFFF7FFF3FFEFFFEDFFEBFFEAFFEBFFECFFEEFFF1FFF5FFF9FFFD",
		INIT_2F=>X"FFF3FFF8FFFD00010006000B000E0012001400150015001500130010000D0009",
		INIT_30=>X"0012000F000A00050000FFFBFFF7FFF2FFEEFFECFFEAFFE9FFE9FFEAFFECFFF0",
		INIT_31=>X"FFE8FFEAFFEDFFF1FFF6FFFB00010006000B000F001300150017001700170015",
		INIT_32=>X"001A001A001800150011000C00070001FFFCFFF6FFF1FFEDFFEAFFE8FFE6FFE6",
		INIT_33=>X"FFE5FFE3FFE3FFE4FFE7FFEAFFEFFFF4FFFA00000006000B001000150018001A",
		INIT_34=>X"0017001B001D001E001D001C00180014000F00090003FFFCFFF6FFF0FFEBFFE8",
		INIT_35=>X"FFEFFFE9FFE4FFE1FFDFFFDFFFE0FFE3FFE6FFECFFF2FFF8FFFF0006000C0012",
		INIT_36=>X"0006000D0014001A001F0022002300230021001D00180012000C0004FFFDFFF6",
		INIT_37=>X"0007FFFEFFF5FFEDFFE6FFE0FFDCFFD9FFD8FFD9FFDCFFE1FFE7FFEEFFF6FFFE",
		INIT_38=>X"FFE8FFF2FFFC0006000F0018001F00250029002B002B00290025001F00180010",
		INIT_39=>X"002900200016000AFFFFFFF4FFE9FFE0FFD9FFD3FFCFFFCEFFD0FFD3FFD8FFE0",
		INIT_3A=>X"FFC3FFCAFFD3FFDFFFEBFFF800060012001E0028002F00350038003800350030",
		INIT_3B=>X"0050004D0046003C002F002100110001FFF2FFE3FFD6FFCCFFC4FFBFFFBDFFBE",
		INIT_3C=>X"FF9AFF97FF99FFA0FFABFFBAFFCBFFDEFFF200060019002A00380044004C0050",
		INIT_3D=>X"007C008A00910091008A007D006B0055003C00210007FFEDFFD5FFC0FFAFFFA2",
		INIT_3E=>X"FF5CFF34FF19FF0BFF09FF13FF27FF42FF64FF8BFFB4FFDD0006002B004C0067",
		INIT_3F=>X"0467044C042003E5039C034702E80282021801AC014100DA007A0022FFD4FF92",
		INIT_40=>X"FEA4FEA5FEC9FF12FF82001600C8019102670341041204D0057105EA06360650",
		INIT_41=>X"FFE10016004C007E00A800C400CF00C600A900780037FFE9FF96FF44FEFBFEC3",
		INIT_42=>X"0065007000720068005300350011FFE9FFC1FF9EFF82FF70FF6CFF76FF8EFFB3",
		INIT_43=>X"0033001D0004FFE9FFD0FFBAFFAAFFA2FFA3FFADFFBFFFD8FFF6001600350050",
		INIT_44=>X"FFD7FFC8FFBEFFBAFFBDFFC6FFD5FFE9FFFF0016002B003D0049004F004D0044",
		INIT_45=>X"FFCCFFD5FFE2FFF20004001600260032003A003D0039003100230011FFFDFFE9",
		INIT_46=>X"000700150022002B00300031002D002400180009FFF9FFE9FFDBFFD1FFCAFFC9",
		INIT_47=>X"002900290024001C00110004FFF6FFEAFFDFFFD7FFD2FFD2FFD7FFDFFFEBFFF9",
		INIT_48=>X"000C0000FFF5FFEAFFE1FFDBFFD8FFD9FFDEFFE6FFF1FFFD000A0015001F0026",
		INIT_49=>X"FFE3FFDEFFDDFFDFFFE4FFECFFF60000000B0015001D002200240023001E0016",
		INIT_4A=>X"FFE9FFF0FFF90003000D0015001B001F0020001E001900110008FFFDFFF3FFEA",
		INIT_4B=>X"000E0015001A001D001D001A0014000D0004FFFBFFF2FFEAFFE4FFE1FFE1FFE3",
		INIT_4C=>X"001A00160011000A0001FFF9FFF1FFEAFFE6FFE4FFE4FFE7FFECFFF4FFFC0005",
		INIT_4D=>X"FFFFFFF7FFF0FFEBFFE7FFE6FFE7FFEAFFF0FFF7FFFF0007000E00140019001A",
		INIT_4E=>X"FFE8FFE8FFE9FFEDFFF3FFF900010008000F00140017001800170013000E0007",
		INIT_4F=>X"FFF5FFFC0003000A000F00140016001700150011000B0004FFFDFFF6FFF0FFEB",
		INIT_50=>X"00100013001500150013000E00090002FFFBFFF5FFEFFFEBFFE9FFE9FFEBFFF0",
		INIT_51=>X"0011000C00070000FFFAFFF4FFEFFFECFFEAFFEBFFEDFFF2FFF7FFFE0004000B",
		INIT_52=>X"FFF8FFF3FFEFFFECFFEBFFECFFEFFFF4FFF900000006000C0010001300140013",
		INIT_53=>X"FFECFFEEFFF1FFF6FFFB00010007000C0010001300130012000F000A0005FFFF",
		INIT_54=>X"FFFD00030008000D0010001200120010000D00080003FFFDFFF7FFF2FFEFFFED",
		INIT_55=>X"001000120011000F000B00070001FFFBFFF6FFF2FFEFFFEDFFEDFFEFFFF3FFF8",
		INIT_56=>X"000A00050000FFFAFFF5FFF1FFEFFFEEFFEEFFF1FFF4FFF9FFFF00040009000E",
		INIT_57=>X"FFF4FFF1FFEFFFEEFFEFFFF2FFF6FFFB00000006000A000E001000110010000E",
		INIT_58=>X"FFF0FFF3FFF7FFFC00020007000B000E00100011000F000C00080003FFFEFFF9",
		INIT_59=>X"00030008000C000F00100010000E000B00070002FFFDFFF8FFF3FFF0FFEFFFEF",
		INIT_5A=>X"0010000F000D000A00050000FFFBFFF7FFF3FFF0FFEFFFEFFFF1FFF5FFF9FFFE",
		INIT_5B=>X"0004FFFFFFFAFFF6FFF2FFF0FFEFFFF0FFF2FFF6FFFAFFFF00040009000D000F",
		INIT_5C=>X"FFF1FFF0FFEFFFF1FFF3FFF7FFFC00010006000A000D000F0010000F000C0009",
		INIT_5D=>X"FFF4FFF8FFFD00020007000B000E000F000F000E000B00070003FFFEFFF9FFF5",
		INIT_5E=>X"0008000C000E000F000F000D000A00060001FFFCFFF8FFF4FFF1FFF0FFF0FFF1",
		INIT_5F=>X"000F000D000900050000FFFBFFF6FFF3FFF0FFF0FFF0FFF2FFF5FFFAFFFE0003",
		INIT_60=>X"FFFEFFFAFFF5FFF2FFF0FFF0FFF0FFF3FFF6FFFB000000050009000D000F0010",
		INIT_61=>X"FFF0FFF0FFF1FFF4FFF8FFFC00010006000A000D000F000F000E000C00080003",
		INIT_62=>X"FFF9FFFE00030007000B000E000F000F000E000B00070002FFFDFFF8FFF4FFF1",
		INIT_63=>X"000C000F0010000F000D000A00060001FFFCFFF7FFF3FFF1FFEFFFF0FFF1FFF5",
		INIT_64=>X"000D00090004FFFFFFFAFFF6FFF2FFF0FFEFFFF0FFF2FFF6FFFAFFFF00040009",
		INIT_65=>X"FFF9FFF5FFF1FFEFFFEFFFF0FFF3FFF7FFFB00000005000A000D000F0010000F",
		INIT_66=>X"FFEFFFF0FFF3FFF8FFFD00020007000B000E00100010000F000C00080003FFFE",
		INIT_67=>X"FFFE00030008000C000F00110010000E000B00070002FFFCFFF7FFF3FFF0FFEF",
		INIT_68=>X"001000110010000E000A00060000FFFBFFF6FFF2FFEFFFEEFFEFFFF1FFF4FFF9",
		INIT_69=>X"00090004FFFFFFF9FFF4FFF1FFEEFFEEFFEFFFF1FFF5FFFA00000005000A000E",
		INIT_6A=>X"FFF3FFEFFFEDFFEDFFEFFFF2FFF6FFFB00010007000B000F001100120010000E",
		INIT_6B=>X"FFEFFFF2FFF7FFFD00030008000D0010001200120010000D00080003FFFDFFF8",
		INIT_6C=>X"0005000A000F0012001300130010000C00070001FFFBFFF6FFF1FFEEFFECFFED",
		INIT_6D=>X"001400130010000C00060000FFF9FFF4FFEFFFECFFEBFFECFFEFFFF3FFF8FFFF",
		INIT_6E=>X"0004FFFEFFF7FFF2FFEDFFEBFFEAFFECFFEFFFF4FFFA00000007000C00110013",
		INIT_6F=>X"FFEBFFE9FFE9FFEBFFEFFFF5FFFB00020009000E00130015001500130010000B",
		INIT_70=>X"FFF0FFF6FFFD0004000B00110015001700160014000F000A0003FFFCFFF5FFF0",
		INIT_71=>X"000E00130017001800170014000F00080001FFF9FFF3FFEDFFE9FFE8FFE8FFEB",
		INIT_72=>X"00190014000E0007FFFFFFF7FFF0FFEAFFE7FFE6FFE7FFEBFFF0FFF7FFFF0007",
		INIT_73=>X"FFFCFFF4FFECFFE7FFE4FFE4FFE6FFEAFFF1FFF90001000A00110016001A001A",
		INIT_74=>X"FFE1FFE1FFE4FFEAFFF2FFFB0004000D0014001A001D001D001A0015000E0005",
		INIT_75=>X"FFF3FFFD000800110019001E0020001F001B0015000D0003FFF9FFF0FFE9FFE3",
		INIT_76=>X"001E002300240022001D0015000B0000FFF6FFECFFE4FFDFFFDDFFDEFFE3FFEA",
		INIT_77=>X"001F0015000AFFFDFFF1FFE6FFDEFFD9FFD8FFDBFFE1FFEAFFF50000000C0016",
		INIT_78=>X"FFEBFFDFFFD7FFD2FFD2FFD7FFDFFFEAFFF600040011001C0024002900290026",
		INIT_79=>X"FFCAFFD1FFDBFFE9FFF9000900180024002D00310030002B002200150007FFF9",
		INIT_7A=>X"FFFD0011002300310039003D003A0032002600160004FFF2FFE2FFD5FFCCFFC9",
		INIT_7B=>X"004D004F0049003D002B0016FFFFFFE9FFD5FFC6FFBDFFBAFFBEFFC8FFD7FFE9",
		INIT_7C=>X"00350016FFF6FFD8FFBFFFADFFA3FFA2FFAAFFBAFFD0FFE90004001D00330044",
		INIT_7D=>X"FF8EFF76FF6CFF70FF82FF9EFFC1FFE900110035005300680072007000650050",
		INIT_7E=>X"FEFBFF44FF96FFE90037007800A900C600CF00C400A8007E004C0016FFE1FFB3",
		INIT_7F=>X"063605EA057104D0041203410267019100C80016FF82FF12FEC9FEA5FEA4FEC3",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_08,
		DOPADOP=>dopadop_08,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_09: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"000FFFFF00000FFFFF00000FFFFFC00003FFFFC00003FFFFC00003FFFFC00000",
		INITP_01=>X"F00000FFFFF00000FFFFFC00003FFFFC00003FFFFC00003FFFFC00000FFFFF00",
		INITP_02=>X"FFFF000003FFFFC00003FFFFC00003FFFFC00003FFFFC00000FFFFF00000FFFF",
		INITP_03=>X"003FFFFC00003FFFFC00003FFFFC00003FFFFF00000FFFFF00000FFFFF00000F",
		INITP_04=>X"C00003FFFFC00003FFFFC00003FFFFF00000FFFFF00000FFFFF00000FFFFF000",
		INITP_05=>X"FFFC00003FFFFC00000FFFFF00000FFFFF00000FFFFF00000FFFFF000003FFFF",
		INITP_06=>X"03FFFFC00000FFFFF00000FFFFF00000FFFFF00000FFFFFC00003FFFFC00003F",
		INITP_07=>X"00000FFFFF00000FFFFF00000FFFFF00000FFFFFC00003FFFFC00003FFFFC000",
		INITP_08=>X"FFF0003FFF0003FFF0000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF0000",
		INITP_09=>X"FFC000FFFC000FFFF0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC0003",
		INITP_0A=>X"FF0003FFF0003FFFC000FFFC000FFFC000FFFF0003FFF0003FFF0003FFFC000F",
		INITP_0B=>X"FC000FFFC0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC000FFFF0003F",
		INITP_0C=>X"F0003FFFC000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF0000FFFC000FF",
		INITP_0D=>X"C000FFFF0003FFF0003FFF0003FFFC000FFFC000FFFC000FFFF0003FFF0003FF",
		INITP_0E=>X"0000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF0003FFFC000FFFC000FFF",
		INITP_0F=>X"0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF",
		INIT_00=>X"FEA4FEA5FEC9FF12FF82001600C8019102670341041204D0057105EA06360650",
		INIT_01=>X"FFE10016004C007E00A800C400CF00C600A900780037FFE9FF96FF44FEFBFEC3",
		INIT_02=>X"0065007000720068005300350011FFE9FFC1FF9EFF82FF70FF6CFF76FF8EFFB3",
		INIT_03=>X"0033001D0004FFE9FFD0FFBAFFAAFFA2FFA3FFADFFBFFFD8FFF6001600350050",
		INIT_04=>X"FFD7FFC8FFBEFFBAFFBDFFC6FFD5FFE9FFFF0016002B003D0049004F004D0044",
		INIT_05=>X"FFCCFFD5FFE2FFF20004001600260032003A003D0039003100230011FFFDFFE9",
		INIT_06=>X"000700150022002B00300031002D002400180009FFF9FFE9FFDBFFD1FFCAFFC9",
		INIT_07=>X"002900290024001C00110004FFF6FFEAFFDFFFD7FFD2FFD2FFD7FFDFFFEBFFF9",
		INIT_08=>X"000C0000FFF5FFEAFFE1FFDBFFD8FFD9FFDEFFE6FFF1FFFD000A0015001F0026",
		INIT_09=>X"FFE3FFDEFFDDFFDFFFE4FFECFFF60000000B0015001D002200240023001E0016",
		INIT_0A=>X"FFE9FFF0FFF90003000D0015001B001F0020001E001900110008FFFDFFF3FFEA",
		INIT_0B=>X"000E0015001A001D001D001A0014000D0004FFFBFFF2FFEAFFE4FFE1FFE1FFE3",
		INIT_0C=>X"001A00160011000A0001FFF9FFF1FFEAFFE6FFE4FFE4FFE7FFECFFF4FFFC0005",
		INIT_0D=>X"FFFFFFF7FFF0FFEBFFE7FFE6FFE7FFEAFFF0FFF7FFFF0007000E00140019001A",
		INIT_0E=>X"FFE8FFE8FFE9FFEDFFF3FFF900010008000F00140017001800170013000E0007",
		INIT_0F=>X"FFF5FFFC0003000A000F00140016001700150011000B0004FFFDFFF6FFF0FFEB",
		INIT_10=>X"00100013001500150013000E00090002FFFBFFF5FFEFFFEBFFE9FFE9FFEBFFF0",
		INIT_11=>X"0011000C00070000FFFAFFF4FFEFFFECFFEAFFEBFFEDFFF2FFF7FFFE0004000B",
		INIT_12=>X"FFF8FFF3FFEFFFECFFEBFFECFFEFFFF4FFF900000006000C0010001300140013",
		INIT_13=>X"FFECFFEEFFF1FFF6FFFB00010007000C0010001300130012000F000A0005FFFF",
		INIT_14=>X"FFFD00030008000D0010001200120010000D00080003FFFDFFF7FFF2FFEFFFED",
		INIT_15=>X"001000120011000F000B00070001FFFBFFF6FFF2FFEFFFEDFFEDFFEFFFF3FFF8",
		INIT_16=>X"000A00050000FFFAFFF5FFF1FFEFFFEEFFEEFFF1FFF4FFF9FFFF00040009000E",
		INIT_17=>X"FFF4FFF1FFEFFFEEFFEFFFF2FFF6FFFB00000006000A000E001000110010000E",
		INIT_18=>X"FFF0FFF3FFF7FFFC00020007000B000E00100011000F000C00080003FFFEFFF9",
		INIT_19=>X"00030008000C000F00100010000E000B00070002FFFDFFF8FFF3FFF0FFEFFFEF",
		INIT_1A=>X"0010000F000D000A00050000FFFBFFF7FFF3FFF0FFEFFFEFFFF1FFF5FFF9FFFE",
		INIT_1B=>X"0004FFFFFFFAFFF6FFF2FFF0FFEFFFF0FFF2FFF6FFFAFFFF00040009000D000F",
		INIT_1C=>X"FFF1FFF0FFEFFFF1FFF3FFF7FFFC00010006000A000D000F0010000F000C0009",
		INIT_1D=>X"FFF4FFF8FFFD00020007000B000E000F000F000E000B00070003FFFEFFF9FFF5",
		INIT_1E=>X"0008000C000E000F000F000D000A00060001FFFCFFF8FFF4FFF1FFF0FFF0FFF1",
		INIT_1F=>X"000F000D000900050000FFFBFFF6FFF3FFF0FFF0FFF0FFF2FFF5FFFAFFFE0003",
		INIT_20=>X"FFFEFFFAFFF5FFF2FFF0FFF0FFF0FFF3FFF6FFFB000000050009000D000F0010",
		INIT_21=>X"FFF0FFF0FFF1FFF4FFF8FFFC00010006000A000D000F000F000E000C00080003",
		INIT_22=>X"FFF9FFFE00030007000B000E000F000F000E000B00070002FFFDFFF8FFF4FFF1",
		INIT_23=>X"000C000F0010000F000D000A00060001FFFCFFF7FFF3FFF1FFEFFFF0FFF1FFF5",
		INIT_24=>X"000D00090004FFFFFFFAFFF6FFF2FFF0FFEFFFF0FFF2FFF6FFFAFFFF00040009",
		INIT_25=>X"FFF9FFF5FFF1FFEFFFEFFFF0FFF3FFF7FFFB00000005000A000D000F0010000F",
		INIT_26=>X"FFEFFFF0FFF3FFF8FFFD00020007000B000E00100010000F000C00080003FFFE",
		INIT_27=>X"FFFE00030008000C000F00110010000E000B00070002FFFCFFF7FFF3FFF0FFEF",
		INIT_28=>X"001000110010000E000A00060000FFFBFFF6FFF2FFEFFFEEFFEFFFF1FFF4FFF9",
		INIT_29=>X"00090004FFFFFFF9FFF4FFF1FFEEFFEEFFEFFFF1FFF5FFFA00000005000A000E",
		INIT_2A=>X"FFF3FFEFFFEDFFEDFFEFFFF2FFF6FFFB00010007000B000F001100120010000E",
		INIT_2B=>X"FFEFFFF2FFF7FFFD00030008000D0010001200120010000D00080003FFFDFFF8",
		INIT_2C=>X"0005000A000F0012001300130010000C00070001FFFBFFF6FFF1FFEEFFECFFED",
		INIT_2D=>X"001400130010000C00060000FFF9FFF4FFEFFFECFFEBFFECFFEFFFF3FFF8FFFF",
		INIT_2E=>X"0004FFFEFFF7FFF2FFEDFFEBFFEAFFECFFEFFFF4FFFA00000007000C00110013",
		INIT_2F=>X"FFEBFFE9FFE9FFEBFFEFFFF5FFFB00020009000E00130015001500130010000B",
		INIT_30=>X"FFF0FFF6FFFD0004000B00110015001700160014000F000A0003FFFCFFF5FFF0",
		INIT_31=>X"000E00130017001800170014000F00080001FFF9FFF3FFEDFFE9FFE8FFE8FFEB",
		INIT_32=>X"00190014000E0007FFFFFFF7FFF0FFEAFFE7FFE6FFE7FFEBFFF0FFF7FFFF0007",
		INIT_33=>X"FFFCFFF4FFECFFE7FFE4FFE4FFE6FFEAFFF1FFF90001000A00110016001A001A",
		INIT_34=>X"FFE1FFE1FFE4FFEAFFF2FFFB0004000D0014001A001D001D001A0015000E0005",
		INIT_35=>X"FFF3FFFD000800110019001E0020001F001B0015000D0003FFF9FFF0FFE9FFE3",
		INIT_36=>X"001E002300240022001D0015000B0000FFF6FFECFFE4FFDFFFDDFFDEFFE3FFEA",
		INIT_37=>X"001F0015000AFFFDFFF1FFE6FFDEFFD9FFD8FFDBFFE1FFEAFFF50000000C0016",
		INIT_38=>X"FFEBFFDFFFD7FFD2FFD2FFD7FFDFFFEAFFF600040011001C0024002900290026",
		INIT_39=>X"FFCAFFD1FFDBFFE9FFF9000900180024002D00310030002B002200150007FFF9",
		INIT_3A=>X"FFFD0011002300310039003D003A0032002600160004FFF2FFE2FFD5FFCCFFC9",
		INIT_3B=>X"004D004F0049003D002B0016FFFFFFE9FFD5FFC6FFBDFFBAFFBEFFC8FFD7FFE9",
		INIT_3C=>X"00350016FFF6FFD8FFBFFFADFFA3FFA2FFAAFFBAFFD0FFE90004001D00330044",
		INIT_3D=>X"FF8EFF76FF6CFF70FF82FF9EFFC1FFE900110035005300680072007000650050",
		INIT_3E=>X"FEFBFF44FF96FFE90037007800A900C600CF00C400A8007E004C0016FFE1FFB3",
		INIT_3F=>X"063605EA057104D0041203410267019100C80016FF82FF12FEC9FEA5FEA4FEC3",
		INIT_40=>X"0065FFCBFF24FE8DFE28FE11FE5DFF15003401A7034F0501069207D508A708F0",
		INIT_41=>X"00900061001CFFCCFF80FF47FF2FFF3DFF73FFCA0034009D00F30121011B00DA",
		INIT_42=>X"006D006E005A00340001FFCCFF9FFF82FF7BFF8FFFB9FFF30033006D009500A2",
		INIT_43=>X"0031004A00550051003C001BFFF4FFCDFFAFFF9FFFA1FFB6FFD9000500320057",
		INIT_44=>X"FFF90016002F00400045003D0029000CFFECFFCFFFBAFFB2FFB9FFCDFFEC0010",
		INIT_45=>X"FFD6FFEA0002001A002E00390039002F001B0001FFE7FFD0FFC3FFC0FFCAFFDE",
		INIT_46=>X"FFD0FFD4FFE0FFF30008001D002C0032003000240010FFFAFFE4FFD2FFC9FFCB",
		INIT_47=>X"FFE0FFD7FFD5FFDBFFE9FFFA000D001E0029002D0027001A0008FFF4FFE2FFD5",
		INIT_48=>X"FFFCFFECFFE0FFDAFFDAFFE2FFF000000011001F00270027002000130001FFF0",
		INIT_49=>X"00140006FFF7FFEAFFE0FFDCFFDFFFE8FFF600050014001F00240022001A000C",
		INIT_4A=>X"001E0019000F0001FFF4FFE8FFE1FFDFFFE4FFEEFFFB000A0016001F0021001D",
		INIT_4B=>X"0018001C001B0014000AFFFDFFF1FFE7FFE2FFE2FFE8FFF30000000D0017001E",
		INIT_4C=>X"000700120019001B001800100005FFF9FFEEFFE7FFE3FFE6FFEDFFF700040010",
		INIT_4D=>X"FFF5FFFF000A0013001800190015000C0002FFF6FFEDFFE7FFE5FFE9FFF1FFFC",
		INIT_4E=>X"FFE9FFEFFFF80003000D00140018001700110009FFFEFFF4FFEBFFE7FFE7FFEC",
		INIT_4F=>X"FFEAFFE9FFECFFF3FFFC0006000F001500170014000E0005FFFBFFF1FFEBFFE8",
		INIT_50=>X"FFF5FFEEFFEAFFEAFFEEFFF6FFFF00080010001500150012000B0002FFF8FFF0",
		INIT_51=>X"0005FFFCFFF3FFEDFFEBFFECFFF1FFF90002000B001100150014000F0008FFFE",
		INIT_52=>X"0010000A0002FFF9FFF1FFEDFFEBFFEEFFF4FFFC0005000D001200140012000D",
		INIT_53=>X"00130012000E0007FFFFFFF7FFF0FFECFFECFFF0FFF6FFFF0007000E00130013",
		INIT_54=>X"000B001000120011000C0004FFFCFFF5FFEFFFEDFFEEFFF2FFF9000100090010",
		INIT_55=>X"FFFF0006000D00110012000F00090002FFFAFFF3FFEEFFEDFFEFFFF5FFFC0004",
		INIT_56=>X"FFF3FFF900010008000E00110011000D0007FFFFFFF8FFF1FFEEFFEEFFF1FFF7",
		INIT_57=>X"FFEEFFF0FFF5FFFC0003000A000F00110010000B0004FFFDFFF6FFF0FFEEFFEF",
		INIT_58=>X"FFF2FFEFFFEFFFF2FFF7FFFE0006000C00100011000E00090002FFFAFFF4FFF0",
		INIT_59=>X"FFFDFFF6FFF1FFEFFFF0FFF3FFF900010008000D00100010000C0007FFFFFFF8",
		INIT_5A=>X"00090002FFFBFFF5FFF0FFEFFFF1FFF5FFFC0003000A000E0010000F000B0004",
		INIT_5B=>X"000F000C00070000FFF9FFF3FFF0FFEFFFF2FFF7FFFE0005000B000F0010000E",
		INIT_5C=>X"000E0010000F000B0004FFFDFFF7FFF2FFEFFFF0FFF4FFF900000007000D0010",
		INIT_5D=>X"0005000B000F0010000D00090002FFFBFFF5FFF1FFEFFFF1FFF5FFFC00030009",
		INIT_5E=>X"FFF900000007000C000F000F000C00070000FFF9FFF3FFF0FFF0FFF2FFF7FFFE",
		INIT_5F=>X"FFF1FFF5FFFB00020009000D000F000E000B0005FFFEFFF7FFF2FFF0FFF0FFF4",
		INIT_60=>X"FFF0FFF0FFF2FFF7FFFE0005000B000E000F000D00090002FFFBFFF5FFF1FFF0",
		INIT_61=>X"FFF7FFF2FFF0FFF0FFF3FFF900000007000C000F000F000C00070000FFF9FFF4",
		INIT_62=>X"0003FFFCFFF5FFF1FFEFFFF1FFF5FFFB00020009000D0010000F000B0005FFFE",
		INIT_63=>X"000D00070000FFF9FFF4FFF0FFEFFFF2FFF7FFFD0004000B000F0010000E0009",
		INIT_64=>X"0010000F000B0005FFFEFFF7FFF2FFEFFFF0FFF3FFF900000007000C000F0010",
		INIT_65=>X"000B000F0010000E000A0003FFFCFFF5FFF1FFEFFFF0FFF5FFFB00020009000E",
		INIT_66=>X"FFFF0007000C00100010000D00080001FFF9FFF3FFF0FFEFFFF1FFF6FFFD0004",
		INIT_67=>X"FFF4FFFA00020009000E00110010000C0006FFFEFFF7FFF2FFEFFFEFFFF2FFF8",
		INIT_68=>X"FFEEFFF0FFF6FFFD0004000B00100011000F000A0003FFFCFFF5FFF0FFEEFFF0",
		INIT_69=>X"FFF1FFEEFFEEFFF1FFF8FFFF0007000D00110011000E00080001FFF9FFF3FFEF",
		INIT_6A=>X"FFFCFFF5FFEFFFEDFFEEFFF3FFFA00020009000F00120011000D0006FFFFFFF7",
		INIT_6B=>X"00090001FFF9FFF2FFEEFFEDFFEFFFF5FFFC0004000C001100120010000B0004",
		INIT_6C=>X"0013000E0007FFFFFFF6FFF0FFECFFECFFF0FFF7FFFF0007000E001200130010",
		INIT_6D=>X"001200140012000D0005FFFCFFF4FFEEFFEBFFEDFFF1FFF90002000A00100013",
		INIT_6E=>X"0008000F001400150011000B0002FFF9FFF1FFECFFEBFFEDFFF3FFFC0005000D",
		INIT_6F=>X"FFF80002000B00120015001500100008FFFFFFF6FFEEFFEAFFEAFFEEFFF5FFFE",
		INIT_70=>X"FFEBFFF1FFFB0005000E001400170015000F0006FFFCFFF3FFECFFE9FFEAFFF0",
		INIT_71=>X"FFE7FFE7FFEBFFF4FFFE00090011001700180014000D0003FFF8FFEFFFE9FFE8",
		INIT_72=>X"FFF1FFE9FFE5FFE7FFEDFFF60002000C0015001900180013000AFFFFFFF5FFEC",
		INIT_73=>X"0004FFF7FFEDFFE6FFE3FFE7FFEEFFF9000500100018001B001900120007FFFC",
		INIT_74=>X"0017000D0000FFF3FFE8FFE2FFE2FFE7FFF1FFFD000A0014001B001C00180010",
		INIT_75=>X"0021001F0016000AFFFBFFEEFFE4FFDFFFE1FFE8FFF40001000F0019001E001E",
		INIT_76=>X"001A00220024001F00140005FFF6FFE8FFDFFFDCFFE0FFEAFFF700060014001D",
		INIT_77=>X"00010013002000270027001F00110000FFF0FFE2FFDAFFDAFFE0FFECFFFC000C",
		INIT_78=>X"FFE2FFF40008001A0027002D0029001E000DFFFAFFE9FFDBFFD5FFD7FFE0FFF0",
		INIT_79=>X"FFC9FFD2FFE4FFFA0010002400300032002C001D0008FFF3FFE0FFD4FFD0FFD5",
		INIT_7A=>X"FFCAFFC0FFC3FFD0FFE70001001B002F00390039002E001A0002FFEAFFD6FFCB",
		INIT_7B=>X"FFECFFCDFFB9FFB2FFBAFFCFFFEC000C0029003D00450040002F0016FFF9FFDE",
		INIT_7C=>X"00320005FFD9FFB6FFA1FF9FFFAFFFCDFFF4001B003C00510055004A00310010",
		INIT_7D=>X"0095006D0033FFF3FFB9FF8FFF7BFF82FF9FFFCC00010034005A006E006D0057",
		INIT_7E=>X"011B012100F3009D0034FFCAFF73FF3DFF2FFF47FF80FFCC001C0061009000A2",
		INIT_7F=>X"08A707D506920501034F01A70034FF15FE5DFE11FE28FE8DFF24FFCB006500DA",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_09,
		DOPADOP=>dopadop_09,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_10: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFF0003FFF0003FFF0000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF0000",
		INITP_01=>X"FFC000FFFC000FFFF0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC0003",
		INITP_02=>X"FF0003FFF0003FFFC000FFFC000FFFC000FFFF0003FFF0003FFF0003FFFC000F",
		INITP_03=>X"FC000FFFC0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC000FFFF0003F",
		INITP_04=>X"F0003FFFC000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF0000FFFC000FF",
		INITP_05=>X"C000FFFF0003FFF0003FFF0003FFFC000FFFC000FFFC000FFFF0003FFF0003FF",
		INITP_06=>X"0000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF0003FFFC000FFFC000FFF",
		INITP_07=>X"0003FFF0003FFF0003FFF0000FFFC000FFFC000FFFC0003FFF0003FFF0003FFF",
		INITP_08=>X"003FF003FFC00FFC00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF000",
		INITP_09=>X"3FF003FF003FF003FF000FFC00FFC00FFC00FFC00FFC00FFF003FF003FF003FF",
		INITP_0A=>X"C003FF003FF003FF003FF003FF003FFC00FFC00FFC00FFC00FFC00FFC003FF00",
		INITP_0B=>X"0FFC00FFC00FFF003FF003FF003FF003FF003FF000FFC00FFC00FFC00FFC00FF",
		INITP_0C=>X"FC00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FFC00FFC00FFC0",
		INITP_0D=>X"03FF000FFC00FFC00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF000F",
		INITP_0E=>X"FF003FF003FF003FFC00FFC00FFC00FFC00FFC00FFC003FF003FF003FF003FF0",
		INITP_0F=>X"003FF003FF003FF003FF003FF000FFC00FFC00FFC00FFC00FFC00FFF003FF003",
		INIT_00=>X"0065FFCBFF24FE8DFE28FE11FE5DFF15003401A7034F0501069207D508A708F0",
		INIT_01=>X"00900061001CFFCCFF80FF47FF2FFF3DFF73FFCA0034009D00F30121011B00DA",
		INIT_02=>X"006D006E005A00340001FFCCFF9FFF82FF7BFF8FFFB9FFF30033006D009500A2",
		INIT_03=>X"0031004A00550051003C001BFFF4FFCDFFAFFF9FFFA1FFB6FFD9000500320057",
		INIT_04=>X"FFF90016002F00400045003D0029000CFFECFFCFFFBAFFB2FFB9FFCDFFEC0010",
		INIT_05=>X"FFD6FFEA0002001A002E00390039002F001B0001FFE7FFD0FFC3FFC0FFCAFFDE",
		INIT_06=>X"FFD0FFD4FFE0FFF30008001D002C0032003000240010FFFAFFE4FFD2FFC9FFCB",
		INIT_07=>X"FFE0FFD7FFD5FFDBFFE9FFFA000D001E0029002D0027001A0008FFF4FFE2FFD5",
		INIT_08=>X"FFFCFFECFFE0FFDAFFDAFFE2FFF000000011001F00270027002000130001FFF0",
		INIT_09=>X"00140006FFF7FFEAFFE0FFDCFFDFFFE8FFF600050014001F00240022001A000C",
		INIT_0A=>X"001E0019000F0001FFF4FFE8FFE1FFDFFFE4FFEEFFFB000A0016001F0021001D",
		INIT_0B=>X"0018001C001B0014000AFFFDFFF1FFE7FFE2FFE2FFE8FFF30000000D0017001E",
		INIT_0C=>X"000700120019001B001800100005FFF9FFEEFFE7FFE3FFE6FFEDFFF700040010",
		INIT_0D=>X"FFF5FFFF000A0013001800190015000C0002FFF6FFEDFFE7FFE5FFE9FFF1FFFC",
		INIT_0E=>X"FFE9FFEFFFF80003000D00140018001700110009FFFEFFF4FFEBFFE7FFE7FFEC",
		INIT_0F=>X"FFEAFFE9FFECFFF3FFFC0006000F001500170014000E0005FFFBFFF1FFEBFFE8",
		INIT_10=>X"FFF5FFEEFFEAFFEAFFEEFFF6FFFF00080010001500150012000B0002FFF8FFF0",
		INIT_11=>X"0005FFFCFFF3FFEDFFEBFFECFFF1FFF90002000B001100150014000F0008FFFE",
		INIT_12=>X"0010000A0002FFF9FFF1FFEDFFEBFFEEFFF4FFFC0005000D001200140012000D",
		INIT_13=>X"00130012000E0007FFFFFFF7FFF0FFECFFECFFF0FFF6FFFF0007000E00130013",
		INIT_14=>X"000B001000120011000C0004FFFCFFF5FFEFFFEDFFEEFFF2FFF9000100090010",
		INIT_15=>X"FFFF0006000D00110012000F00090002FFFAFFF3FFEEFFEDFFEFFFF5FFFC0004",
		INIT_16=>X"FFF3FFF900010008000E00110011000D0007FFFFFFF8FFF1FFEEFFEEFFF1FFF7",
		INIT_17=>X"FFEEFFF0FFF5FFFC0003000A000F00110010000B0004FFFDFFF6FFF0FFEEFFEF",
		INIT_18=>X"FFF2FFEFFFEFFFF2FFF7FFFE0006000C00100011000E00090002FFFAFFF4FFF0",
		INIT_19=>X"FFFDFFF6FFF1FFEFFFF0FFF3FFF900010008000D00100010000C0007FFFFFFF8",
		INIT_1A=>X"00090002FFFBFFF5FFF0FFEFFFF1FFF5FFFC0003000A000E0010000F000B0004",
		INIT_1B=>X"000F000C00070000FFF9FFF3FFF0FFEFFFF2FFF7FFFE0005000B000F0010000E",
		INIT_1C=>X"000E0010000F000B0004FFFDFFF7FFF2FFEFFFF0FFF4FFF900000007000D0010",
		INIT_1D=>X"0005000B000F0010000D00090002FFFBFFF5FFF1FFEFFFF1FFF5FFFC00030009",
		INIT_1E=>X"FFF900000007000C000F000F000C00070000FFF9FFF3FFF0FFF0FFF2FFF7FFFE",
		INIT_1F=>X"FFF1FFF5FFFB00020009000D000F000E000B0005FFFEFFF7FFF2FFF0FFF0FFF4",
		INIT_20=>X"FFF0FFF0FFF2FFF7FFFE0005000B000E000F000D00090002FFFBFFF5FFF1FFF0",
		INIT_21=>X"FFF7FFF2FFF0FFF0FFF3FFF900000007000C000F000F000C00070000FFF9FFF4",
		INIT_22=>X"0003FFFCFFF5FFF1FFEFFFF1FFF5FFFB00020009000D0010000F000B0005FFFE",
		INIT_23=>X"000D00070000FFF9FFF4FFF0FFEFFFF2FFF7FFFD0004000B000F0010000E0009",
		INIT_24=>X"0010000F000B0005FFFEFFF7FFF2FFEFFFF0FFF3FFF900000007000C000F0010",
		INIT_25=>X"000B000F0010000E000A0003FFFCFFF5FFF1FFEFFFF0FFF5FFFB00020009000E",
		INIT_26=>X"FFFF0007000C00100010000D00080001FFF9FFF3FFF0FFEFFFF1FFF6FFFD0004",
		INIT_27=>X"FFF4FFFA00020009000E00110010000C0006FFFEFFF7FFF2FFEFFFEFFFF2FFF8",
		INIT_28=>X"FFEEFFF0FFF6FFFD0004000B00100011000F000A0003FFFCFFF5FFF0FFEEFFF0",
		INIT_29=>X"FFF1FFEEFFEEFFF1FFF8FFFF0007000D00110011000E00080001FFF9FFF3FFEF",
		INIT_2A=>X"FFFCFFF5FFEFFFEDFFEEFFF3FFFA00020009000F00120011000D0006FFFFFFF7",
		INIT_2B=>X"00090001FFF9FFF2FFEEFFEDFFEFFFF5FFFC0004000C001100120010000B0004",
		INIT_2C=>X"0013000E0007FFFFFFF6FFF0FFECFFECFFF0FFF7FFFF0007000E001200130010",
		INIT_2D=>X"001200140012000D0005FFFCFFF4FFEEFFEBFFEDFFF1FFF90002000A00100013",
		INIT_2E=>X"0008000F001400150011000B0002FFF9FFF1FFECFFEBFFEDFFF3FFFC0005000D",
		INIT_2F=>X"FFF80002000B00120015001500100008FFFFFFF6FFEEFFEAFFEAFFEEFFF5FFFE",
		INIT_30=>X"FFEBFFF1FFFB0005000E001400170015000F0006FFFCFFF3FFECFFE9FFEAFFF0",
		INIT_31=>X"FFE7FFE7FFEBFFF4FFFE00090011001700180014000D0003FFF8FFEFFFE9FFE8",
		INIT_32=>X"FFF1FFE9FFE5FFE7FFEDFFF60002000C0015001900180013000AFFFFFFF5FFEC",
		INIT_33=>X"0004FFF7FFEDFFE6FFE3FFE7FFEEFFF9000500100018001B001900120007FFFC",
		INIT_34=>X"0017000D0000FFF3FFE8FFE2FFE2FFE7FFF1FFFD000A0014001B001C00180010",
		INIT_35=>X"0021001F0016000AFFFBFFEEFFE4FFDFFFE1FFE8FFF40001000F0019001E001E",
		INIT_36=>X"001A00220024001F00140005FFF6FFE8FFDFFFDCFFE0FFEAFFF700060014001D",
		INIT_37=>X"00010013002000270027001F00110000FFF0FFE2FFDAFFDAFFE0FFECFFFC000C",
		INIT_38=>X"FFE2FFF40008001A0027002D0029001E000DFFFAFFE9FFDBFFD5FFD7FFE0FFF0",
		INIT_39=>X"FFC9FFD2FFE4FFFA0010002400300032002C001D0008FFF3FFE0FFD4FFD0FFD5",
		INIT_3A=>X"FFCAFFC0FFC3FFD0FFE70001001B002F00390039002E001A0002FFEAFFD6FFCB",
		INIT_3B=>X"FFECFFCDFFB9FFB2FFBAFFCFFFEC000C0029003D00450040002F0016FFF9FFDE",
		INIT_3C=>X"00320005FFD9FFB6FFA1FF9FFFAFFFCDFFF4001B003C00510055004A00310010",
		INIT_3D=>X"0095006D0033FFF3FFB9FF8FFF7BFF82FF9FFFCC00010034005A006E006D0057",
		INIT_3E=>X"011B012100F3009D0034FFCAFF73FF3DFF2FFF47FF80FFCC001C0061009000A2",
		INIT_3F=>X"08A707D506920501034F01A70034FF15FE5DFE11FE28FE8DFF24FFCB006500DA",
		INIT_40=>X"003C0109018B018600E3FFC3FE7CFD83FD50FE33003C032E0687099C0BC80C90",
		INIT_41=>X"002CFFC4FF6BFF45FF63FFBF003C00AB00E200C7005CFFC3FF31FEDFFEF4FF74",
		INIT_42=>X"FFB7FFF5003A006C007700560013FFC5FF89FF77FF98FFE1003B0083009D007E",
		INIT_43=>X"004C002BFFF8FFC7FFA9FFABFFCC00020038005C005E003C0003FFC6FF9CFF96",
		INIT_44=>X"FFBDFFC8FFE7001100350046003D001DFFF1FFC9FFB4FFBBFFDC000B00370050",
		INIT_45=>X"003100370028000AFFE7FFCDFFC4FFD2FFF100160033003E00320013FFEBFFCB",
		INIT_46=>X"FFE2FFD1FFD1FFE3FFFF001C002F003100200003FFE4FFCFFFCBFFDBFFF90019",
		INIT_47=>X"0009001F002A00250012FFF8FFE0FFD4FFD7FFE90004001E002D002B0019FFFD",
		INIT_48=>X"0008FFF1FFDFFFD9FFE1FFF5000D002000270020000DFFF4FFDFFFD6FFDCFFF0",
		INIT_49=>X"FFEBFFFE00120020002100170003FFEEFFDFFFDCFFE6FFFA001000200024001B",
		INIT_4A=>X"001B000EFFFBFFEAFFE0FFE2FFEF00020014001F001E0012FFFFFFECFFDFFFDF",
		INIT_4B=>X"FFE3FFE8FFF700080017001D0018000AFFF8FFE9FFE1FFE5FFF300050016001E",
		INIT_4C=>X"0018001A00120003FFF3FFE7FFE4FFEBFFFA000B0018001C00150007FFF5FFE8",
		INIT_4D=>X"FFEFFFE7FFE8FFF20001000F00180018000F0000FFF1FFE7FFE6FFEEFFFD000D",
		INIT_4E=>X"00060012001800140009FFFAFFEDFFE7FFEAFFF50003001100180016000CFFFD",
		INIT_4F=>X"0003FFF6FFECFFE9FFEEFFFA00080013001700120006FFF8FFECFFE8FFECFFF7",
		INIT_50=>X"FFF30000000C00140015000D0001FFF4FFEBFFEAFFF1FFFD000A001400160010",
		INIT_51=>X"00120008FFFCFFF1FFEBFFEDFFF60002000E00140013000BFFFEFFF2FFEBFFEB",
		INIT_52=>X"FFECFFF0FFFA00070010001400100006FFFAFFEFFFEBFFEEFFF80004000F0014",
		INIT_53=>X"00120012000C0001FFF6FFEEFFECFFF2FFFD000800110013000E0003FFF8FFEE",
		INIT_54=>X"FFF3FFEDFFEEFFF60001000C00120011000AFFFFFFF4FFEDFFEDFFF4FFFF000A",
		INIT_55=>X"0005000E0012000F0006FFFBFFF1FFEDFFF0FFF80003000D001200100008FFFD",
		INIT_56=>X"0002FFF7FFF0FFEEFFF3FFFC0007000F0011000D0004FFF9FFF0FFEDFFF1FFFA",
		INIT_57=>X"FFF60000000A00100010000A0000FFF5FFEFFFEFFFF4FFFE000900100011000B",
		INIT_58=>X"000E0006FFFCFFF3FFEFFFF1FFF80002000C0010000F0008FFFEFFF4FFEFFFF0",
		INIT_59=>X"FFEFFFF3FFFC0006000E0010000D0004FFFAFFF2FFEFFFF2FFFA0004000D0010",
		INIT_5A=>X"000F000F000A0000FFF6FFF0FFEFFFF5FFFE0008000F0010000B0002FFF8FFF1",
		INIT_5B=>X"FFF4FFEFFFF1FFF80002000B0010000E0008FFFEFFF5FFF0FFF0FFF600000009",
		INIT_5C=>X"0005000D0010000C0004FFFBFFF2FFEFFFF2FFFA0004000C0010000E0006FFFC",
		INIT_5D=>X"0001FFF7FFF1FFF0FFF5FFFD0007000E000F000B0003FFF9FFF2FFEFFFF3FFFC",
		INIT_5E=>X"FFF80001000A000F000E0008FFFFFFF6FFF0FFF0FFF6FFFF0009000F000F000A",
		INIT_5F=>X"000D0005FFFBFFF3FFF0FFF2FFF90003000B000F000E0007FFFDFFF4FFF0FFF1",
		INIT_60=>X"FFF0FFF4FFFD0007000E000F000B0003FFF9FFF2FFF0FFF3FFFB0005000D0010",
		INIT_61=>X"000F000F0009FFFFFFF6FFF0FFF0FFF6FFFF0008000E000F000A0001FFF8FFF1",
		INIT_62=>X"FFF3FFEFFFF2FFF90003000B000F000E0007FFFDFFF5FFF0FFF1FFF70001000A",
		INIT_63=>X"0006000E0010000C0004FFFAFFF2FFEFFFF2FFFB0004000C0010000D0005FFFC",
		INIT_64=>X"0000FFF6FFF0FFF0FFF5FFFE0008000E0010000B0002FFF8FFF1FFEFFFF4FFFC",
		INIT_65=>X"FFF80002000B0010000F0008FFFEFFF5FFEFFFF0FFF60000000A000F000F0009",
		INIT_66=>X"000D0004FFFAFFF2FFEFFFF2FFFA0004000D0010000E0006FFFCFFF3FFEFFFF1",
		INIT_67=>X"FFEFFFF4FFFE0008000F0010000C0002FFF8FFF1FFEFFFF3FFFC0006000E0010",
		INIT_68=>X"001100100009FFFEFFF4FFEFFFEFFFF50000000A00100010000A0000FFF6FFF0",
		INIT_69=>X"FFF1FFEDFFF0FFF90004000D0011000F0007FFFCFFF3FFEEFFF0FFF70002000B",
		INIT_6A=>X"000800100012000D0003FFF8FFF0FFEDFFF1FFFB0006000F0012000E0005FFFA",
		INIT_6B=>X"FFFFFFF4FFEDFFEDFFF4FFFF000A00110012000C0001FFF6FFEEFFEDFFF3FFFD",
		INIT_6C=>X"FFF80003000E001300110008FFFDFFF2FFECFFEEFFF60001000C00120012000A",
		INIT_6D=>X"000F0004FFF8FFEEFFEBFFEFFFFA00060010001400100007FFFAFFF0FFECFFEE",
		INIT_6E=>X"FFEBFFF2FFFE000B00130014000E0002FFF6FFEDFFEBFFF1FFFC000800120014",
		INIT_6F=>X"00160014000AFFFDFFF1FFEAFFEBFFF40001000D00150014000C0000FFF3FFEB",
		INIT_70=>X"FFECFFE8FFECFFF800060012001700130008FFFAFFEEFFE9FFECFFF600030010",
		INIT_71=>X"000C0016001800110003FFF5FFEAFFE7FFEDFFFA00090014001800120006FFF7",
		INIT_72=>X"FFFDFFEEFFE6FFE7FFF10000000F00180018000F0001FFF2FFE8FFE7FFEFFFFD",
		INIT_73=>X"FFF500070015001C0018000BFFFAFFEBFFE4FFE7FFF300030012001A0018000D",
		INIT_74=>X"00160005FFF3FFE5FFE1FFE9FFF8000A0018001D00170008FFF7FFE8FFE3FFE8",
		INIT_75=>X"FFDFFFECFFFF0012001E001F00140002FFEFFFE2FFE0FFEAFFFB000E001B001E",
		INIT_76=>X"002400200010FFFAFFE6FFDCFFDFFFEE00030017002100200012FFFEFFEBFFDF",
		INIT_77=>X"FFDCFFD6FFDFFFF4000D002000270020000DFFF5FFE1FFD9FFDFFFF10008001B",
		INIT_78=>X"0019002B002D001E0004FFE9FFD7FFD4FFE0FFF800120025002A001F0009FFF0",
		INIT_79=>X"FFF9FFDBFFCBFFCFFFE4000300200031002F001CFFFFFFE3FFD1FFD1FFE2FFFD",
		INIT_7A=>X"FFEB00130032003E00330016FFF1FFD2FFC4FFCDFFE7000A0028003700310019",
		INIT_7B=>X"0037000BFFDCFFBBFFB4FFC9FFF1001D003D004600350011FFE7FFC8FFBDFFCB",
		INIT_7C=>X"FF9CFFC60003003C005E005C00380002FFCCFFABFFA9FFC7FFF8002B004C0050",
		INIT_7D=>X"009D0083003BFFE1FF98FF77FF89FFC5001300560077006C003AFFF5FFB7FF96",
		INIT_7E=>X"FEF4FEDFFF31FFC3005C00C700E200AB003CFFBFFF63FF45FF6BFFC4002C007E",
		INIT_7F=>X"0BC8099C0687032E003CFE33FD50FD83FE7CFFC300E30186018B0109003CFF74",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_10,
		DOPADOP=>dopadop_10,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_11: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"003FF003FFC00FFC00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF000",
		INITP_01=>X"3FF003FF003FF003FF000FFC00FFC00FFC00FFC00FFC00FFF003FF003FF003FF",
		INITP_02=>X"C003FF003FF003FF003FF003FF003FFC00FFC00FFC00FFC00FFC00FFC003FF00",
		INITP_03=>X"0FFC00FFC00FFF003FF003FF003FF003FF003FF000FFC00FFC00FFC00FFC00FF",
		INITP_04=>X"FC00FFC00FFC00FFC00FFC003FF003FF003FF003FF003FF003FFC00FFC00FFC0",
		INITP_05=>X"03FF000FFC00FFC00FFC00FFC00FFC00FFF003FF003FF003FF003FF003FF000F",
		INITP_06=>X"FF003FF003FF003FFC00FFC00FFC00FFC00FFC00FFC003FF003FF003FF003FF0",
		INITP_07=>X"003FF003FF003FF003FF003FF000FFC00FFC00FFC00FFC00FFC00FFF003FF003",
		INITP_08=>X"00FC03FC0FF03FC03F00FF03FC03F00FF03FC0FF00FC03FC0FF00FC03FC0FF00",
		INITP_09=>X"FF00FC03FC0FF00FC03F00FF03FC03F00FF03FC03F00FF03FC0FF00FC03FC0FF",
		INITP_0A=>X"C03F00FC03FC0FF00FC03FC0FF00FC03F00FF03FC03F00FF03FC03F00FC03FC0",
		INITP_0B=>X"3FC03F00FF03FC0FF00FC03FC0FF00FC03FC0FF03FC03F00FF03FC03F00FF03F",
		INITP_0C=>X"F03FC03F00FF03FC03F00FF03FC0FF00FC03FC0FF00FC03FC0FF03FC03F00FF0",
		INITP_0D=>X"0FF00FC03F00FF03FC03F00FF03FC03F00FC03FC0FF00FC03FC0FF00FC03F00F",
		INITP_0E=>X"FC0FF00FC03FC0FF03FC03F00FF03FC03F00FF03FC03F00FC03FC0FF00FC03FC",
		INITP_0F=>X"03FC0FF00FC03FC0FF00FC03FC0FF03FC03F00FF03FC03F00FF03FC0FF00FC03",
		INIT_00=>X"003C0109018B018600E3FFC3FE7CFD83FD50FE33003C032E0687099C0BC80C90",
		INIT_01=>X"002CFFC4FF6BFF45FF63FFBF003C00AB00E200C7005CFFC3FF31FEDFFEF4FF74",
		INIT_02=>X"FFB7FFF5003A006C007700560013FFC5FF89FF77FF98FFE1003B0083009D007E",
		INIT_03=>X"004C002BFFF8FFC7FFA9FFABFFCC00020038005C005E003C0003FFC6FF9CFF96",
		INIT_04=>X"FFBDFFC8FFE7001100350046003D001DFFF1FFC9FFB4FFBBFFDC000B00370050",
		INIT_05=>X"003100370028000AFFE7FFCDFFC4FFD2FFF100160033003E00320013FFEBFFCB",
		INIT_06=>X"FFE2FFD1FFD1FFE3FFFF001C002F003100200003FFE4FFCFFFCBFFDBFFF90019",
		INIT_07=>X"0009001F002A00250012FFF8FFE0FFD4FFD7FFE90004001E002D002B0019FFFD",
		INIT_08=>X"0008FFF1FFDFFFD9FFE1FFF5000D002000270020000DFFF4FFDFFFD6FFDCFFF0",
		INIT_09=>X"FFEBFFFE00120020002100170003FFEEFFDFFFDCFFE6FFFA001000200024001B",
		INIT_0A=>X"001B000EFFFBFFEAFFE0FFE2FFEF00020014001F001E0012FFFFFFECFFDFFFDF",
		INIT_0B=>X"FFE3FFE8FFF700080017001D0018000AFFF8FFE9FFE1FFE5FFF300050016001E",
		INIT_0C=>X"0018001A00120003FFF3FFE7FFE4FFEBFFFA000B0018001C00150007FFF5FFE8",
		INIT_0D=>X"FFEFFFE7FFE8FFF20001000F00180018000F0000FFF1FFE7FFE6FFEEFFFD000D",
		INIT_0E=>X"00060012001800140009FFFAFFEDFFE7FFEAFFF50003001100180016000CFFFD",
		INIT_0F=>X"0003FFF6FFECFFE9FFEEFFFA00080013001700120006FFF8FFECFFE8FFECFFF7",
		INIT_10=>X"FFF30000000C00140015000D0001FFF4FFEBFFEAFFF1FFFD000A001400160010",
		INIT_11=>X"00120008FFFCFFF1FFEBFFEDFFF60002000E00140013000BFFFEFFF2FFEBFFEB",
		INIT_12=>X"FFECFFF0FFFA00070010001400100006FFFAFFEFFFEBFFEEFFF80004000F0014",
		INIT_13=>X"00120012000C0001FFF6FFEEFFECFFF2FFFD000800110013000E0003FFF8FFEE",
		INIT_14=>X"FFF3FFEDFFEEFFF60001000C00120011000AFFFFFFF4FFEDFFEDFFF4FFFF000A",
		INIT_15=>X"0005000E0012000F0006FFFBFFF1FFEDFFF0FFF80003000D001200100008FFFD",
		INIT_16=>X"0002FFF7FFF0FFEEFFF3FFFC0007000F0011000D0004FFF9FFF0FFEDFFF1FFFA",
		INIT_17=>X"FFF60000000A00100010000A0000FFF5FFEFFFEFFFF4FFFE000900100011000B",
		INIT_18=>X"000E0006FFFCFFF3FFEFFFF1FFF80002000C0010000F0008FFFEFFF4FFEFFFF0",
		INIT_19=>X"FFEFFFF3FFFC0006000E0010000D0004FFFAFFF2FFEFFFF2FFFA0004000D0010",
		INIT_1A=>X"000F000F000A0000FFF6FFF0FFEFFFF5FFFE0008000F0010000B0002FFF8FFF1",
		INIT_1B=>X"FFF4FFEFFFF1FFF80002000B0010000E0008FFFEFFF5FFF0FFF0FFF600000009",
		INIT_1C=>X"0005000D0010000C0004FFFBFFF2FFEFFFF2FFFA0004000C0010000E0006FFFC",
		INIT_1D=>X"0001FFF7FFF1FFF0FFF5FFFD0007000E000F000B0003FFF9FFF2FFEFFFF3FFFC",
		INIT_1E=>X"FFF80001000A000F000E0008FFFFFFF6FFF0FFF0FFF6FFFF0009000F000F000A",
		INIT_1F=>X"000D0005FFFBFFF3FFF0FFF2FFF90003000B000F000E0007FFFDFFF4FFF0FFF1",
		INIT_20=>X"FFF0FFF4FFFD0007000E000F000B0003FFF9FFF2FFF0FFF3FFFB0005000D0010",
		INIT_21=>X"000F000F0009FFFFFFF6FFF0FFF0FFF6FFFF0008000E000F000A0001FFF8FFF1",
		INIT_22=>X"FFF3FFEFFFF2FFF90003000B000F000E0007FFFDFFF5FFF0FFF1FFF70001000A",
		INIT_23=>X"0006000E0010000C0004FFFAFFF2FFEFFFF2FFFB0004000C0010000D0005FFFC",
		INIT_24=>X"0000FFF6FFF0FFF0FFF5FFFE0008000E0010000B0002FFF8FFF1FFEFFFF4FFFC",
		INIT_25=>X"FFF80002000B0010000F0008FFFEFFF5FFEFFFF0FFF60000000A000F000F0009",
		INIT_26=>X"000D0004FFFAFFF2FFEFFFF2FFFA0004000D0010000E0006FFFCFFF3FFEFFFF1",
		INIT_27=>X"FFEFFFF4FFFE0008000F0010000C0002FFF8FFF1FFEFFFF3FFFC0006000E0010",
		INIT_28=>X"001100100009FFFEFFF4FFEFFFEFFFF50000000A00100010000A0000FFF6FFF0",
		INIT_29=>X"FFF1FFEDFFF0FFF90004000D0011000F0007FFFCFFF3FFEEFFF0FFF70002000B",
		INIT_2A=>X"000800100012000D0003FFF8FFF0FFEDFFF1FFFB0006000F0012000E0005FFFA",
		INIT_2B=>X"FFFFFFF4FFEDFFEDFFF4FFFF000A00110012000C0001FFF6FFEEFFEDFFF3FFFD",
		INIT_2C=>X"FFF80003000E001300110008FFFDFFF2FFECFFEEFFF60001000C00120012000A",
		INIT_2D=>X"000F0004FFF8FFEEFFEBFFEFFFFA00060010001400100007FFFAFFF0FFECFFEE",
		INIT_2E=>X"FFEBFFF2FFFE000B00130014000E0002FFF6FFEDFFEBFFF1FFFC000800120014",
		INIT_2F=>X"00160014000AFFFDFFF1FFEAFFEBFFF40001000D00150014000C0000FFF3FFEB",
		INIT_30=>X"FFECFFE8FFECFFF800060012001700130008FFFAFFEEFFE9FFECFFF600030010",
		INIT_31=>X"000C0016001800110003FFF5FFEAFFE7FFEDFFFA00090014001800120006FFF7",
		INIT_32=>X"FFFDFFEEFFE6FFE7FFF10000000F00180018000F0001FFF2FFE8FFE7FFEFFFFD",
		INIT_33=>X"FFF500070015001C0018000BFFFAFFEBFFE4FFE7FFF300030012001A0018000D",
		INIT_34=>X"00160005FFF3FFE5FFE1FFE9FFF8000A0018001D00170008FFF7FFE8FFE3FFE8",
		INIT_35=>X"FFDFFFECFFFF0012001E001F00140002FFEFFFE2FFE0FFEAFFFB000E001B001E",
		INIT_36=>X"002400200010FFFAFFE6FFDCFFDFFFEE00030017002100200012FFFEFFEBFFDF",
		INIT_37=>X"FFDCFFD6FFDFFFF4000D002000270020000DFFF5FFE1FFD9FFDFFFF10008001B",
		INIT_38=>X"0019002B002D001E0004FFE9FFD7FFD4FFE0FFF800120025002A001F0009FFF0",
		INIT_39=>X"FFF9FFDBFFCBFFCFFFE4000300200031002F001CFFFFFFE3FFD1FFD1FFE2FFFD",
		INIT_3A=>X"FFEB00130032003E00330016FFF1FFD2FFC4FFCDFFE7000A0028003700310019",
		INIT_3B=>X"0037000BFFDCFFBBFFB4FFC9FFF1001D003D004600350011FFE7FFC8FFBDFFCB",
		INIT_3C=>X"FF9CFFC60003003C005E005C00380002FFCCFFABFFA9FFC7FFF8002B004C0050",
		INIT_3D=>X"009D0083003BFFE1FF98FF77FF89FFC5001300560077006C003AFFF5FFB7FF96",
		INIT_3E=>X"FEF4FEDFFF31FFC3005C00C700E200AB003CFFBFFF63FF45FF6BFFC4002C007E",
		INIT_3F=>X"0BC8099C0687032E003CFE33FD50FD83FE7CFFC300E30186018B0109003CFF74",
		INIT_40=>X"007CFF4EFE77FEA6FFE4017702400177FF48FCF5FC40FE7603940A100F771190",
		INIT_41=>X"00A80074FFE8FF63FF46FFAD005800D100BC001BFF57FEFBFF550036010A0133",
		INIT_42=>X"002300690067001BFFB8FF83FFA50009006B00860041FFCAFF72FF7BFFE40067",
		INIT_43=>X"FFBEFFFC003E00560032FFE8FFACFFAAFFE400340061004BFFFEFFAFFF96FFC7",
		INIT_44=>X"FFC7FFBFFFE4001E0043003A0007FFCDFFB6FFD2000F00430049001BFFD8FFAF",
		INIT_45=>X"000CFFDEFFC7FFD70005002F0039001AFFE8FFC5FFCBFFF600290040002AFFF6",
		INIT_46=>X"002F001AFFF2FFD3FFD2FFF2001B00320026FFFEFFD7FFCBFFE5001100320030",
		INIT_47=>X"0013002900220003FFE1FFD4FFE500090027002A000EFFE8FFD2FFDBFFFE0023",
		INIT_48=>X"FFE60003001F00250010FFF0FFDAFFDEFFFA001A0028001AFFF9FFDCFFD8FFF0",
		INIT_49=>X"FFE0FFE1FFF7001300220019FFFEFFE3FFDCFFEE000C002200200007FFE9FFDA",
		INIT_4A=>X"0002FFE9FFE0FFED0007001C001D000AFFEFFFDFFFE6FFFF001900210012FFF6",
		INIT_4B=>X"001B000CFFF3FFE3FFE7FFFC0013001D0012FFFAFFE5FFE3FFF4000E001E0018",
		INIT_4C=>X"000F001A0013FFFEFFEAFFE5FFF2000A001A00180005FFEEFFE3FFEC00030017",
		INIT_4D=>X"FFF10006001600170007FFF2FFE6FFEC000000130019000DFFF7FFE7FFE8FFF9",
		INIT_4E=>X"FFE8FFECFFFD00100018000FFFFBFFEAFFE8FFF7000B001800130001FFEDFFE6",
		INIT_4F=>X"FFFEFFEDFFE9FFF50008001500130003FFF1FFE8FFF00003001300160009FFF5",
		INIT_50=>X"00130006FFF4FFEAFFEF000000100015000BFFF8FFEBFFECFFFA000D00160010",
		INIT_51=>X"000E0014000CFFFBFFEDFFECFFF8000A001400100000FFF0FFEAFFF300050013",
		INIT_52=>X"FFF70007001300110003FFF2FFEBFFF20003001100130008FFF6FFECFFEFFFFD",
		INIT_53=>X"FFECFFF10000000F00130009FFF9FFEDFFEEFFFB000B0013000DFFFEFFEFFFEC",
		INIT_54=>X"FFFBFFEFFFEEFFF900090012000E0000FFF1FFEDFFF50005001100110005FFF5",
		INIT_55=>X"000F0002FFF3FFEDFFF40003000F00110006FFF7FFEEFFF0FFFE000D0012000B",
		INIT_56=>X"000E00110008FFF9FFEFFFF0FFFC000B0011000CFFFEFFF1FFEEFFF800070011",
		INIT_57=>X"FFFA00090011000D0000FFF2FFEEFFF600050010000F0004FFF5FFEEFFF30000",
		INIT_58=>X"FFEEFFF50003000E00100006FFF7FFEFFFF2FFFE000C0011000AFFFBFFF0FFF0",
		INIT_59=>X"FFF9FFF0FFF1FFFC000A0010000BFFFDFFF1FFEFFFF800070010000E0002FFF4",
		INIT_5A=>X"000CFFFFFFF3FFEFFFF70005000F000E0003FFF6FFEFFFF40001000D00100007",
		INIT_5B=>X"000E000F0005FFF8FFEFFFF3FFFF000B00100009FFFBFFF1FFF0FFFB00080010",
		INIT_5C=>X"FFFD000A0010000AFFFDFFF2FFF0FFF90006000F000D0001FFF4FFEFFFF50003",
		INIT_5D=>X"FFF0FFF70005000E000E0003FFF6FFEFFFF40001000D000F0007FFF9FFF0FFF2",
		INIT_5E=>X"FFF8FFF0FFF3FFFF000B000F0008FFFBFFF1FFF1FFFB0008000F000BFFFFFFF3",
		INIT_5F=>X"000AFFFDFFF2FFF0FFF90007000F000D0001FFF4FFF0FFF60003000E000E0005",
		INIT_60=>X"000E000E0003FFF6FFF0FFF40001000D000F0007FFF9FFF0FFF2FFFD000A0010",
		INIT_61=>X"FFFF000B000F0008FFFBFFF1FFF1FFFB0008000F000BFFFFFFF3FFF0FFF80005",
		INIT_62=>X"FFF0FFF90007000F000D0001FFF4FFEFFFF60003000E000E0005FFF7FFF0FFF3",
		INIT_63=>X"FFF5FFEFFFF40001000D000F0006FFF9FFF0FFF2FFFD000A0010000AFFFDFFF2",
		INIT_64=>X"0008FFFBFFF0FFF1FFFB00090010000BFFFFFFF3FFEFFFF80005000F000E0003",
		INIT_65=>X"0010000D0001FFF4FFEFFFF60003000E000F0005FFF7FFEFFFF3FFFF000C0010",
		INIT_66=>X"0002000E00100007FFF8FFEFFFF1FFFD000B0010000AFFFCFFF1FFF0FFF90007",
		INIT_67=>X"FFF0FFFB000A0011000CFFFEFFF2FFEFFFF700060010000E0003FFF5FFEEFFF4",
		INIT_68=>X"FFF3FFEEFFF50004000F00100005FFF6FFEEFFF20000000D00110009FFFAFFF0",
		INIT_69=>X"0007FFF8FFEEFFF1FFFE000C0011000BFFFCFFF0FFEFFFF900080011000E0000",
		INIT_6A=>X"0012000DFFFEFFF0FFEEFFF700060011000F0003FFF4FFEDFFF30002000F0011",
		INIT_6B=>X"0005001100110005FFF5FFEDFFF10000000E00120009FFF9FFEEFFEFFFFB000B",
		INIT_6C=>X"FFEFFFFE000D0013000BFFFBFFEEFFEDFFF900090013000F0000FFF1FFECFFF5",
		INIT_6D=>X"FFEFFFECFFF60008001300110003FFF2FFEBFFF20003001100130007FFF7FFEC",
		INIT_6E=>X"0005FFF3FFEAFFF0000000100014000AFFF8FFECFFEDFFFB000C0014000EFFFD",
		INIT_6F=>X"0016000DFFFAFFECFFEBFFF8000B001500100000FFEFFFEAFFF4000600130013",
		INIT_70=>X"0009001600130003FFF0FFE8FFF10003001300150008FFF5FFE9FFEDFFFE0010",
		INIT_71=>X"FFED000100130018000BFFF7FFE8FFEAFFFB000F00180010FFFDFFECFFE8FFF5",
		INIT_72=>X"FFE8FFE7FFF7000D001900130000FFECFFE6FFF20007001700160006FFF1FFE6",
		INIT_73=>X"0003FFECFFE3FFEE00050018001A000AFFF2FFE5FFEAFFFE0013001A000FFFF9",
		INIT_74=>X"001E000EFFF4FFE3FFE5FFFA0012001D0013FFFCFFE7FFE3FFF3000C001B0017",
		INIT_75=>X"001200210019FFFFFFE6FFDFFFEF000A001D001C0007FFEDFFE0FFE900020018",
		INIT_76=>X"FFE9000700200022000CFFEEFFDCFFE3FFFE001900220013FFF7FFE1FFE0FFF6",
		INIT_77=>X"FFD8FFDCFFF9001A0028001AFFFAFFDEFFDAFFF000100025001F0003FFE6FFDA",
		INIT_78=>X"FFFEFFDBFFD2FFE8000E002A00270009FFE5FFD4FFE10003002200290013FFF0",
		INIT_79=>X"00320011FFE5FFCBFFD7FFFE00260032001BFFF2FFD2FFD3FFF2001A002F0023",
		INIT_7A=>X"002A00400029FFF6FFCBFFC5FFE8001A0039002F0005FFD7FFC7FFDE000C0030",
		INIT_7B=>X"FFD8001B00490043000FFFD2FFB6FFCD0007003A0043001EFFE4FFBFFFC7FFF6",
		INIT_7C=>X"FF96FFAFFFFE004B00610034FFE4FFAAFFACFFE800320056003EFFFCFFBEFFAF",
		INIT_7D=>X"FFE4FF7BFF72FFCA00410086006B0009FFA5FF83FFB8001B006700690023FFC7",
		INIT_7E=>X"010A0036FF55FEFBFF57001B00BC00D10058FFADFF46FF63FFE8007400A80067",
		INIT_7F=>X"0F770A100394FE76FC40FCF5FF48017702400177FFE4FEA6FE77FF4E007C0133",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_11,
		DOPADOP=>dopadop_11,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_12: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"00FC03FC0FF03FC03F00FF03FC03F00FF03FC0FF00FC03FC0FF00FC03FC0FF00",
		INITP_01=>X"FF00FC03FC0FF00FC03F00FF03FC03F00FF03FC03F00FF03FC0FF00FC03FC0FF",
		INITP_02=>X"C03F00FC03FC0FF00FC03FC0FF00FC03F00FF03FC03F00FF03FC03F00FC03FC0",
		INITP_03=>X"3FC03F00FF03FC0FF00FC03FC0FF00FC03FC0FF03FC03F00FF03FC03F00FF03F",
		INITP_04=>X"F03FC03F00FF03FC03F00FF03FC0FF00FC03FC0FF00FC03FC0FF03FC03F00FF0",
		INITP_05=>X"0FF00FC03F00FF03FC03F00FF03FC03F00FC03FC0FF00FC03FC0FF00FC03F00F",
		INITP_06=>X"FC0FF00FC03FC0FF03FC03F00FF03FC03F00FF03FC03F00FC03FC0FF00FC03FC",
		INITP_07=>X"03FC0FF00FC03FC0FF00FC03FC0FF03FC03F00FF03FC03F00FF03FC0FF00FC03",
		INITP_08=>X"03F0FC3F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC0",
		INITP_09=>X"3F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F",
		INITP_0A=>X"F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC",
		INITP_0B=>X"C3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0",
		INITP_0C=>X"0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0F",
		INITP_0D=>X"FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3F03C",
		INITP_0E=>X"C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3F03C0F03F0",
		INITP_0F=>X"0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3F03C0F03F0FC3F03",
		INIT_00=>X"007CFF4EFE77FEA6FFE4017702400177FF48FCF5FC40FE7603940A100F771190",
		INIT_01=>X"00A80074FFE8FF63FF46FFAD005800D100BC001BFF57FEFBFF550036010A0133",
		INIT_02=>X"002300690067001BFFB8FF83FFA50009006B00860041FFCAFF72FF7BFFE40067",
		INIT_03=>X"FFBEFFFC003E00560032FFE8FFACFFAAFFE400340061004BFFFEFFAFFF96FFC7",
		INIT_04=>X"FFC7FFBFFFE4001E0043003A0007FFCDFFB6FFD2000F00430049001BFFD8FFAF",
		INIT_05=>X"000CFFDEFFC7FFD70005002F0039001AFFE8FFC5FFCBFFF600290040002AFFF6",
		INIT_06=>X"002F001AFFF2FFD3FFD2FFF2001B00320026FFFEFFD7FFCBFFE5001100320030",
		INIT_07=>X"0013002900220003FFE1FFD4FFE500090027002A000EFFE8FFD2FFDBFFFE0023",
		INIT_08=>X"FFE60003001F00250010FFF0FFDAFFDEFFFA001A0028001AFFF9FFDCFFD8FFF0",
		INIT_09=>X"FFE0FFE1FFF7001300220019FFFEFFE3FFDCFFEE000C002200200007FFE9FFDA",
		INIT_0A=>X"0002FFE9FFE0FFED0007001C001D000AFFEFFFDFFFE6FFFF001900210012FFF6",
		INIT_0B=>X"001B000CFFF3FFE3FFE7FFFC0013001D0012FFFAFFE5FFE3FFF4000E001E0018",
		INIT_0C=>X"000F001A0013FFFEFFEAFFE5FFF2000A001A00180005FFEEFFE3FFEC00030017",
		INIT_0D=>X"FFF10006001600170007FFF2FFE6FFEC000000130019000DFFF7FFE7FFE8FFF9",
		INIT_0E=>X"FFE8FFECFFFD00100018000FFFFBFFEAFFE8FFF7000B001800130001FFEDFFE6",
		INIT_0F=>X"FFFEFFEDFFE9FFF50008001500130003FFF1FFE8FFF00003001300160009FFF5",
		INIT_10=>X"00130006FFF4FFEAFFEF000000100015000BFFF8FFEBFFECFFFA000D00160010",
		INIT_11=>X"000E0014000CFFFBFFEDFFECFFF8000A001400100000FFF0FFEAFFF300050013",
		INIT_12=>X"FFF70007001300110003FFF2FFEBFFF20003001100130008FFF6FFECFFEFFFFD",
		INIT_13=>X"FFECFFF10000000F00130009FFF9FFEDFFEEFFFB000B0013000DFFFEFFEFFFEC",
		INIT_14=>X"FFFBFFEFFFEEFFF900090012000E0000FFF1FFEDFFF50005001100110005FFF5",
		INIT_15=>X"000F0002FFF3FFEDFFF40003000F00110006FFF7FFEEFFF0FFFE000D0012000B",
		INIT_16=>X"000E00110008FFF9FFEFFFF0FFFC000B0011000CFFFEFFF1FFEEFFF800070011",
		INIT_17=>X"FFFA00090011000D0000FFF2FFEEFFF600050010000F0004FFF5FFEEFFF30000",
		INIT_18=>X"FFEEFFF50003000E00100006FFF7FFEFFFF2FFFE000C0011000AFFFBFFF0FFF0",
		INIT_19=>X"FFF9FFF0FFF1FFFC000A0010000BFFFDFFF1FFEFFFF800070010000E0002FFF4",
		INIT_1A=>X"000CFFFFFFF3FFEFFFF70005000F000E0003FFF6FFEFFFF40001000D00100007",
		INIT_1B=>X"000E000F0005FFF8FFEFFFF3FFFF000B00100009FFFBFFF1FFF0FFFB00080010",
		INIT_1C=>X"FFFD000A0010000AFFFDFFF2FFF0FFF90006000F000D0001FFF4FFEFFFF50003",
		INIT_1D=>X"FFF0FFF70005000E000E0003FFF6FFEFFFF40001000D000F0007FFF9FFF0FFF2",
		INIT_1E=>X"FFF8FFF0FFF3FFFF000B000F0008FFFBFFF1FFF1FFFB0008000F000BFFFFFFF3",
		INIT_1F=>X"000AFFFDFFF2FFF0FFF90007000F000D0001FFF4FFF0FFF60003000E000E0005",
		INIT_20=>X"000E000E0003FFF6FFF0FFF40001000D000F0007FFF9FFF0FFF2FFFD000A0010",
		INIT_21=>X"FFFF000B000F0008FFFBFFF1FFF1FFFB0008000F000BFFFFFFF3FFF0FFF80005",
		INIT_22=>X"FFF0FFF90007000F000D0001FFF4FFEFFFF60003000E000E0005FFF7FFF0FFF3",
		INIT_23=>X"FFF5FFEFFFF40001000D000F0006FFF9FFF0FFF2FFFD000A0010000AFFFDFFF2",
		INIT_24=>X"0008FFFBFFF0FFF1FFFB00090010000BFFFFFFF3FFEFFFF80005000F000E0003",
		INIT_25=>X"0010000D0001FFF4FFEFFFF60003000E000F0005FFF7FFEFFFF3FFFF000C0010",
		INIT_26=>X"0002000E00100007FFF8FFEFFFF1FFFD000B0010000AFFFCFFF1FFF0FFF90007",
		INIT_27=>X"FFF0FFFB000A0011000CFFFEFFF2FFEFFFF700060010000E0003FFF5FFEEFFF4",
		INIT_28=>X"FFF3FFEEFFF50004000F00100005FFF6FFEEFFF20000000D00110009FFFAFFF0",
		INIT_29=>X"0007FFF8FFEEFFF1FFFE000C0011000BFFFCFFF0FFEFFFF900080011000E0000",
		INIT_2A=>X"0012000DFFFEFFF0FFEEFFF700060011000F0003FFF4FFEDFFF30002000F0011",
		INIT_2B=>X"0005001100110005FFF5FFEDFFF10000000E00120009FFF9FFEEFFEFFFFB000B",
		INIT_2C=>X"FFEFFFFE000D0013000BFFFBFFEEFFEDFFF900090013000F0000FFF1FFECFFF5",
		INIT_2D=>X"FFEFFFECFFF60008001300110003FFF2FFEBFFF20003001100130007FFF7FFEC",
		INIT_2E=>X"0005FFF3FFEAFFF0000000100014000AFFF8FFECFFEDFFFB000C0014000EFFFD",
		INIT_2F=>X"0016000DFFFAFFECFFEBFFF8000B001500100000FFEFFFEAFFF4000600130013",
		INIT_30=>X"0009001600130003FFF0FFE8FFF10003001300150008FFF5FFE9FFEDFFFE0010",
		INIT_31=>X"FFED000100130018000BFFF7FFE8FFEAFFFB000F00180010FFFDFFECFFE8FFF5",
		INIT_32=>X"FFE8FFE7FFF7000D001900130000FFECFFE6FFF20007001700160006FFF1FFE6",
		INIT_33=>X"0003FFECFFE3FFEE00050018001A000AFFF2FFE5FFEAFFFE0013001A000FFFF9",
		INIT_34=>X"001E000EFFF4FFE3FFE5FFFA0012001D0013FFFCFFE7FFE3FFF3000C001B0017",
		INIT_35=>X"001200210019FFFFFFE6FFDFFFEF000A001D001C0007FFEDFFE0FFE900020018",
		INIT_36=>X"FFE9000700200022000CFFEEFFDCFFE3FFFE001900220013FFF7FFE1FFE0FFF6",
		INIT_37=>X"FFD8FFDCFFF9001A0028001AFFFAFFDEFFDAFFF000100025001F0003FFE6FFDA",
		INIT_38=>X"FFFEFFDBFFD2FFE8000E002A00270009FFE5FFD4FFE10003002200290013FFF0",
		INIT_39=>X"00320011FFE5FFCBFFD7FFFE00260032001BFFF2FFD2FFD3FFF2001A002F0023",
		INIT_3A=>X"002A00400029FFF6FFCBFFC5FFE8001A0039002F0005FFD7FFC7FFDE000C0030",
		INIT_3B=>X"FFD8001B00490043000FFFD2FFB6FFCD0007003A0043001EFFE4FFBFFFC7FFF6",
		INIT_3C=>X"FF96FFAFFFFE004B00610034FFE4FFAAFFACFFE800320056003EFFFCFFBEFFAF",
		INIT_3D=>X"FFE4FF7BFF72FFCA00410086006B0009FFA5FF83FFB8001B006700690023FFC7",
		INIT_3E=>X"010A0036FF55FEFBFF57001B00BC00D10058FFADFF46FF63FFE8007400A80067",
		INIT_3F=>X"0F770A100394FE76FC40FCF5FF48017702400177FFE4FEA6FE77FF4E007C0133",
		INIT_40=>X"FF27FE9DFFED018F0148FF1EFDBEFF52025A02D5FF18FAF4FCC706B3131218B0",
		INIT_41=>X"FFE9FF56FF9C006D00BA0012FF44FF62005800ED004DFF34FF140033012D00A7",
		INIT_42=>X"002CFFAEFF97000A00750049FFBAFF80FFED0078006AFFCDFF6AFFC90076008F",
		INIT_43=>X"0043FFE9FFAAFFD9003D0053FFFCFFA7FFC4003100610012FFA8FFAD0020006C",
		INIT_44=>X"00420012FFC8FFC5000F00460022FFD0FFBAFFFF00470033FFDBFFB1FFED0044",
		INIT_45=>X"00310028FFEAFFC6FFED002D0033FFF5FFC4FFE00026003B0003FFC5FFD2001C",
		INIT_46=>X"001A002F0007FFD4FFDA001100320012FFD9FFD200060033001DFFE0FFCBFFFA",
		INIT_47=>X"00010028001BFFEAFFD5FFF700250023FFF2FFD2FFED00200029FFFCFFD2FFE3",
		INIT_48=>X"FFED001800230000FFDBFFE6001200270009FFDEFFDF000A00280012FFE3FFD9",
		INIT_49=>X"FFE2000500210012FFEAFFDEFFFD00200019FFF0FFDBFFF5001D001FFFF8FFDA",
		INIT_4A=>X"FFE0FFF40017001CFFFCFFE0FFED0012001F0003FFE2FFE7000C0021000AFFE5",
		INIT_4B=>X"FFE7FFE80008001D000CFFEAFFE40002001C0012FFEFFFE2FFFB001A0017FFF5",
		INIT_4C=>X"FFF3FFE5FFF900160016FFF9FFE4FFF300120019FFFFFFE5FFED000E001C0005",
		INIT_4D=>X"0001FFE8FFEE000A00190007FFEBFFEA00050019000CFFEEFFE6FFFF00180012",
		INIT_4E=>X"000DFFF2FFE8FFFD00150011FFF6FFE7FFF700120015FFFCFFE7FFF2000F0018",
		INIT_4F=>X"0014FFFEFFEAFFF2000C00160003FFEBFFEE000700170008FFEEFFEA00020017",
		INIT_50=>X"00150009FFF1FFEB00000014000EFFF5FFEAFFFB00120011FFF9FFE9FFF60010",
		INIT_51=>X"00100011FFFBFFEBFFF5000D00130000FFECFFF1000900150005FFEEFFEE0005",
		INIT_52=>X"000700140006FFF0FFEE00030013000AFFF3FFECFFFE0012000EFFF7FFEBFFF9",
		INIT_53=>X"FFFC0010000EFFF9FFECFFF8000E0011FFFDFFECFFF4000B00130002FFEEFFF1",
		INIT_54=>X"FFF3000900120003FFF0FFF0000500120007FFF2FFEE00010012000BFFF5FFED",
		INIT_55=>X"FFEEFFFF0010000CFFF7FFEDFFFB000F000FFFFBFFEDFFF7000C0011FFFFFFEE",
		INIT_56=>X"FFEEFFF6000A00110001FFEFFFF3000700110005FFF1FFF0000300110009FFF4",
		INIT_57=>X"FFF3FFF000010010000AFFF6FFEFFFFD000F000DFFF9FFEEFFFA000D000FFFFD",
		INIT_58=>X"FFFBFFEFFFF8000B000FFFFFFFEFFFF5000800100002FFF1FFF2000500110006",
		INIT_59=>X"0004FFF2FFF2000300100007FFF4FFF00000000F000BFFF7FFEFFFFC000E000D",
		INIT_5A=>X"000BFFF9FFEFFFFB000D000EFFFCFFEFFFF7000A000F0000FFF0FFF400070010",
		INIT_5B=>X"000F0002FFF1FFF3000500100005FFF3FFF1000200100008FFF6FFF0FFFE000E",
		INIT_5C=>X"000F000AFFF7FFF0FFFD000D000CFFFAFFEFFFF9000B000EFFFEFFF0FFF60009",
		INIT_5D=>X"000A000FFFFFFFF0FFF50007000F0003FFF2FFF2000400100006FFF4FFF10000",
		INIT_5E=>X"0002000F0008FFF5FFF0FFFF000E000BFFF9FFF0FFFB000D000DFFFCFFF0FFF8",
		INIT_5F=>X"FFFA000C000EFFFDFFF0FFF70009000F0001FFF1FFF40006000F0004FFF3FFF2",
		INIT_60=>X"FFF30004000F0006FFF4FFF10001000F0009FFF7FFF0FFFD000E000CFFFAFFF0",
		INIT_61=>X"FFF0FFFC000D000DFFFBFFF0FFF9000B000EFFFFFFF0FFF50008000F0002FFF2",
		INIT_62=>X"FFF1FFF4000600100004FFF2FFF20003000F0007FFF5FFF0FFFF000F000AFFF8",
		INIT_63=>X"FFF6FFF0FFFE000E000BFFF9FFEFFFFA000C000DFFFDFFF0FFF7000A000F0000",
		INIT_64=>X"FFFEFFF0FFF6000800100002FFF1FFF3000500100005FFF3FFF10002000F0009",
		INIT_65=>X"0007FFF4FFF00000000F000AFFF7FFEFFFFC000E000DFFFBFFEFFFF9000B000E",
		INIT_66=>X"000EFFFCFFEFFFF7000B000F0000FFF0FFF4000700100003FFF2FFF200040010",
		INIT_67=>X"00110005FFF2FFF1000200100008FFF5FFEFFFFF000F000BFFF8FFEFFFFB000D",
		INIT_68=>X"000F000DFFFAFFEEFFF9000D000FFFFDFFEFFFF6000A00100001FFF0FFF30006",
		INIT_69=>X"000900110003FFF0FFF1000500110007FFF3FFEF00010011000AFFF6FFEEFFFD",
		INIT_6A=>X"FFFF0011000CFFF7FFEDFFFB000F000FFFFBFFEDFFF7000C0010FFFFFFEEFFF4",
		INIT_6B=>X"FFF5000B00120001FFEEFFF2000700120005FFF0FFF0000300120009FFF3FFEE",
		INIT_6C=>X"FFEE00020013000BFFF4FFECFFFD0011000EFFF8FFECFFF9000E0010FFFCFFED",
		INIT_6D=>X"FFEBFFF7000E0012FFFEFFECFFF3000A00130003FFEEFFF0000600140007FFF1",
		INIT_6E=>X"FFEEFFEE000500150009FFF1FFEC00000013000DFFF5FFEBFFFB00110010FFF9",
		INIT_6F=>X"FFF6FFE9FFF900110012FFFBFFEAFFF5000E00140000FFEBFFF1000900150005",
		INIT_70=>X"0002FFEAFFEE000800170007FFEEFFEB00030016000CFFF2FFEAFFFE00140010",
		INIT_71=>X"000FFFF2FFE7FFFC00150012FFF7FFE7FFF600110015FFFDFFE8FFF2000D0017",
		INIT_72=>X"0018FFFFFFE6FFEE000C00190005FFEAFFEB00070019000AFFEEFFE800010018",
		INIT_73=>X"001C000EFFEDFFE5FFFF00190012FFF3FFE4FFF900160016FFF9FFE5FFF30012",
		INIT_74=>X"0017001AFFFBFFE2FFEF0012001C0002FFE4FFEA000C001D0008FFE8FFE70005",
		INIT_75=>X"000A0021000CFFE7FFE20003001F0012FFEDFFE0FFFC001C0017FFF4FFE0FFF5",
		INIT_76=>X"FFF8001F001DFFF5FFDBFFF000190020FFFDFFDEFFEA001200210005FFE2FFE5",
		INIT_77=>X"FFE300120028000AFFDFFFDE000900270012FFE6FFDB000000230018FFEDFFDA",
		INIT_78=>X"FFD2FFFC00290020FFEDFFD2FFF200230025FFF7FFD5FFEA001B00280001FFD9",
		INIT_79=>X"FFCBFFE0001D00330006FFD2FFD9001200320011FFDAFFD40007002F001AFFE3",
		INIT_7A=>X"FFD2FFC50003003B0026FFE0FFC4FFF50033002DFFEDFFC6FFEA00280031FFFA",
		INIT_7B=>X"FFEDFFB1FFDB00330047FFFFFFBAFFD000220046000FFFC5FFC800120042001C",
		INIT_7C=>X"0020FFADFFA8001200610031FFC4FFA7FFFC0053003DFFD9FFAAFFE900430044",
		INIT_7D=>X"0076FFC9FF6AFFCD006A0078FFEDFF80FFBA00490075000AFF97FFAE002C006C",
		INIT_7E=>X"012D0033FF14FF34004D00ED0058FF62FF44001200BA006DFF9CFF56FFE9008F",
		INIT_7F=>X"131206B3FCC7FAF4FF1802D5025AFF52FDBEFF1E0148018FFFEDFE9DFF2700A7",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_12,
		DOPADOP=>dopadop_12,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_13: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"03F0FC3F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC0",
		INITP_01=>X"3F03C0F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F",
		INITP_02=>X"F03F0FC3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC",
		INITP_03=>X"C3F03C0F03F0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC0F03C0F03F0FC3F03C0",
		INITP_04=>X"0F03F0FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0F",
		INITP_05=>X"FC3F03C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3F03C",
		INITP_06=>X"C0F03C0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3F03C0F03F0",
		INITP_07=>X"0FC3F0FC0F03C0FC3F0FC0F03C0FC3F0FC3F03C0F03F0FC3F03C0F03F0FC3F03",
		INITP_08=>X"0C3C3C3CF0F0F0C3C3C30F0F0F3C3C3C30F0F0F3C3C3CF0F0F0C3C3C3CF0F0F0",
		INITP_09=>X"F0F3C3C3CF0F0F0C3C3C3CF0F0F0C3C3C30F0F0F3C3C3C30F0F0F3C3C3CF0F0F",
		INITP_0A=>X"0F0F3C3C3C30F0F0F3C3C3CF0F0F0C3C3C3CF0F0F0C3C3C30F0F0F3C3C3C30F0",
		INITP_0B=>X"F0F0F0C3C3C30F0F0F3C3C3C30F0F0F3C3C3CF0F0F0C3C3C3CF0F0F0C3C3C30F",
		INITP_0C=>X"C30F0F0C3C3C3CF0F0F0C3C3C3CF0F0F3C3C3C30F0F0F3C3C3C30F0F0C3C3C3C",
		INITP_0D=>X"3C30F0F0F3C3C3C30F0F0C3C3C3CF0F0F0C3C3C3CF0F0F3C3C3C30F0F0F3C3C3",
		INITP_0E=>X"C3C3CF0F0F3C3C3C30F0F0F3C3C3C30F0F0C3C3C3CF0F0F0C3C3C3CF0F0F3C3C",
		INITP_0F=>X"3C3C3CF0F0F0C3C3C3CF0F0F3C3C3C30F0F0F3C3C3C30F0F0C3C3C3CF0F0F0C3",
		INIT_00=>X"FF27FE9DFFED018F0148FF1EFDBEFF52025A02D5FF18FAF4FCC706B3131218B0",
		INIT_01=>X"FFE9FF56FF9C006D00BA0012FF44FF62005800ED004DFF34FF140033012D00A7",
		INIT_02=>X"002CFFAEFF97000A00750049FFBAFF80FFED0078006AFFCDFF6AFFC90076008F",
		INIT_03=>X"0043FFE9FFAAFFD9003D0053FFFCFFA7FFC4003100610012FFA8FFAD0020006C",
		INIT_04=>X"00420012FFC8FFC5000F00460022FFD0FFBAFFFF00470033FFDBFFB1FFED0044",
		INIT_05=>X"00310028FFEAFFC6FFED002D0033FFF5FFC4FFE00026003B0003FFC5FFD2001C",
		INIT_06=>X"001A002F0007FFD4FFDA001100320012FFD9FFD200060033001DFFE0FFCBFFFA",
		INIT_07=>X"00010028001BFFEAFFD5FFF700250023FFF2FFD2FFED00200029FFFCFFD2FFE3",
		INIT_08=>X"FFED001800230000FFDBFFE6001200270009FFDEFFDF000A00280012FFE3FFD9",
		INIT_09=>X"FFE2000500210012FFEAFFDEFFFD00200019FFF0FFDBFFF5001D001FFFF8FFDA",
		INIT_0A=>X"FFE0FFF40017001CFFFCFFE0FFED0012001F0003FFE2FFE7000C0021000AFFE5",
		INIT_0B=>X"FFE7FFE80008001D000CFFEAFFE40002001C0012FFEFFFE2FFFB001A0017FFF5",
		INIT_0C=>X"FFF3FFE5FFF900160016FFF9FFE4FFF300120019FFFFFFE5FFED000E001C0005",
		INIT_0D=>X"0001FFE8FFEE000A00190007FFEBFFEA00050019000CFFEEFFE6FFFF00180012",
		INIT_0E=>X"000DFFF2FFE8FFFD00150011FFF6FFE7FFF700120015FFFCFFE7FFF2000F0018",
		INIT_0F=>X"0014FFFEFFEAFFF2000C00160003FFEBFFEE000700170008FFEEFFEA00020017",
		INIT_10=>X"00150009FFF1FFEB00000014000EFFF5FFEAFFFB00120011FFF9FFE9FFF60010",
		INIT_11=>X"00100011FFFBFFEBFFF5000D00130000FFECFFF1000900150005FFEEFFEE0005",
		INIT_12=>X"000700140006FFF0FFEE00030013000AFFF3FFECFFFE0012000EFFF7FFEBFFF9",
		INIT_13=>X"FFFC0010000EFFF9FFECFFF8000E0011FFFDFFECFFF4000B00130002FFEEFFF1",
		INIT_14=>X"FFF3000900120003FFF0FFF0000500120007FFF2FFEE00010012000BFFF5FFED",
		INIT_15=>X"FFEEFFFF0010000CFFF7FFEDFFFB000F000FFFFBFFEDFFF7000C0011FFFFFFEE",
		INIT_16=>X"FFEEFFF6000A00110001FFEFFFF3000700110005FFF1FFF0000300110009FFF4",
		INIT_17=>X"FFF3FFF000010010000AFFF6FFEFFFFD000F000DFFF9FFEEFFFA000D000FFFFD",
		INIT_18=>X"FFFBFFEFFFF8000B000FFFFFFFEFFFF5000800100002FFF1FFF2000500110006",
		INIT_19=>X"0004FFF2FFF2000300100007FFF4FFF00000000F000BFFF7FFEFFFFC000E000D",
		INIT_1A=>X"000BFFF9FFEFFFFB000D000EFFFCFFEFFFF7000A000F0000FFF0FFF400070010",
		INIT_1B=>X"000F0002FFF1FFF3000500100005FFF3FFF1000200100008FFF6FFF0FFFE000E",
		INIT_1C=>X"000F000AFFF7FFF0FFFD000D000CFFFAFFEFFFF9000B000EFFFEFFF0FFF60009",
		INIT_1D=>X"000A000FFFFFFFF0FFF50007000F0003FFF2FFF2000400100006FFF4FFF10000",
		INIT_1E=>X"0002000F0008FFF5FFF0FFFF000E000BFFF9FFF0FFFB000D000DFFFCFFF0FFF8",
		INIT_1F=>X"FFFA000C000EFFFDFFF0FFF70009000F0001FFF1FFF40006000F0004FFF3FFF2",
		INIT_20=>X"FFF30004000F0006FFF4FFF10001000F0009FFF7FFF0FFFD000E000CFFFAFFF0",
		INIT_21=>X"FFF0FFFC000D000DFFFBFFF0FFF9000B000EFFFFFFF0FFF50008000F0002FFF2",
		INIT_22=>X"FFF1FFF4000600100004FFF2FFF20003000F0007FFF5FFF0FFFF000F000AFFF8",
		INIT_23=>X"FFF6FFF0FFFE000E000BFFF9FFEFFFFA000C000DFFFDFFF0FFF7000A000F0000",
		INIT_24=>X"FFFEFFF0FFF6000800100002FFF1FFF3000500100005FFF3FFF10002000F0009",
		INIT_25=>X"0007FFF4FFF00000000F000AFFF7FFEFFFFC000E000DFFFBFFEFFFF9000B000E",
		INIT_26=>X"000EFFFCFFEFFFF7000B000F0000FFF0FFF4000700100003FFF2FFF200040010",
		INIT_27=>X"00110005FFF2FFF1000200100008FFF5FFEFFFFF000F000BFFF8FFEFFFFB000D",
		INIT_28=>X"000F000DFFFAFFEEFFF9000D000FFFFDFFEFFFF6000A00100001FFF0FFF30006",
		INIT_29=>X"000900110003FFF0FFF1000500110007FFF3FFEF00010011000AFFF6FFEEFFFD",
		INIT_2A=>X"FFFF0011000CFFF7FFEDFFFB000F000FFFFBFFEDFFF7000C0010FFFFFFEEFFF4",
		INIT_2B=>X"FFF5000B00120001FFEEFFF2000700120005FFF0FFF0000300120009FFF3FFEE",
		INIT_2C=>X"FFEE00020013000BFFF4FFECFFFD0011000EFFF8FFECFFF9000E0010FFFCFFED",
		INIT_2D=>X"FFEBFFF7000E0012FFFEFFECFFF3000A00130003FFEEFFF0000600140007FFF1",
		INIT_2E=>X"FFEEFFEE000500150009FFF1FFEC00000013000DFFF5FFEBFFFB00110010FFF9",
		INIT_2F=>X"FFF6FFE9FFF900110012FFFBFFEAFFF5000E00140000FFEBFFF1000900150005",
		INIT_30=>X"0002FFEAFFEE000800170007FFEEFFEB00030016000CFFF2FFEAFFFE00140010",
		INIT_31=>X"000FFFF2FFE7FFFC00150012FFF7FFE7FFF600110015FFFDFFE8FFF2000D0017",
		INIT_32=>X"0018FFFFFFE6FFEE000C00190005FFEAFFEB00070019000AFFEEFFE800010018",
		INIT_33=>X"001C000EFFEDFFE5FFFF00190012FFF3FFE4FFF900160016FFF9FFE5FFF30012",
		INIT_34=>X"0017001AFFFBFFE2FFEF0012001C0002FFE4FFEA000C001D0008FFE8FFE70005",
		INIT_35=>X"000A0021000CFFE7FFE20003001F0012FFEDFFE0FFFC001C0017FFF4FFE0FFF5",
		INIT_36=>X"FFF8001F001DFFF5FFDBFFF000190020FFFDFFDEFFEA001200210005FFE2FFE5",
		INIT_37=>X"FFE300120028000AFFDFFFDE000900270012FFE6FFDB000000230018FFEDFFDA",
		INIT_38=>X"FFD2FFFC00290020FFEDFFD2FFF200230025FFF7FFD5FFEA001B00280001FFD9",
		INIT_39=>X"FFCBFFE0001D00330006FFD2FFD9001200320011FFDAFFD40007002F001AFFE3",
		INIT_3A=>X"FFD2FFC50003003B0026FFE0FFC4FFF50033002DFFEDFFC6FFEA00280031FFFA",
		INIT_3B=>X"FFEDFFB1FFDB00330047FFFFFFBAFFD000220046000FFFC5FFC800120042001C",
		INIT_3C=>X"0020FFADFFA8001200610031FFC4FFA7FFFC0053003DFFD9FFAAFFE900430044",
		INIT_3D=>X"0076FFC9FF6AFFCD006A0078FFEDFF80FFBA00490075000AFF97FFAE002C006C",
		INIT_3E=>X"012D0033FF14FF34004D00ED0058FF62FF44001200BA006DFF9CFF56FFE9008F",
		INIT_3F=>X"131206B3FCC7FAF4FF1802D5025AFF52FDBEFF1E0148018FFFEDFE9DFF2700A7",
		INIT_40=>X"006CFE92FFE601B1FFA7FE0F00F60226FE25FDAC034B0274F9AFFD7614352290",
		INIT_41=>X"007A0066FF62FFBA00BB0019FF2F001A00DBFFA9FF25009800C8FF21FF5B0126",
		INIT_42=>X"FF980036005EFFAFFFB100680036FF83FFE60089FFF7FF71002D008BFFABFF81",
		INIT_43=>X"0005FFAB000F0053FFDAFFB3003A0040FFB3FFD0005B0019FF9AFFFF006AFFE5",
		INIT_44=>X"003A0019FFBDFFF60046FFF7FFBA001A0041FFD4FFC8003B002AFFB8FFE60050",
		INIT_45=>X"FFD200260024FFCFFFE60037000BFFC40003003CFFEDFFC600210031FFD1FFD8",
		INIT_46=>X"FFF7FFD100140029FFE0FFDD00280019FFD0FFF200330000FFCA000C0032FFE6",
		INIT_47=>X"00280005FFD50004002AFFF0FFD900190021FFDDFFE70029000EFFD2FFFC002F",
		INIT_48=>X"FFE7001F0010FFDBFFF80026FFFEFFD9000B0024FFEAFFE0001D0018FFDBFFF0",
		INIT_49=>X"FFF2FFE200150018FFE4FFEE00200009FFDCFFFF0024FFF7FFDD0011001EFFE6",
		INIT_4A=>X"001FFFFCFFE1000B001CFFEDFFE800180012FFE2FFF500200002FFDE00050020",
		INIT_4B=>X"FFF3001B0006FFE20001001DFFF7FFE4000F0017FFEAFFED001A000BFFE2FFFB",
		INIT_4C=>X"FFEFFFEC0015000DFFE6FFF8001B0000FFE40006001AFFF2FFE800130012FFE8",
		INIT_4D=>X"0018FFF7FFE9000E0013FFECFFF100170008FFE6FFFD001AFFFBFFE6000A0017",
		INIT_4E=>X"FFFA0017FFFFFFE800060016FFF3FFEC0011000FFFEAFFF600170003FFE60002",
		INIT_4F=>X"FFEEFFF400140006FFE9FFFF0017FFFAFFEA000A0013FFF0FFF00013000AFFE9",
		INIT_50=>X"0013FFF3FFEF0010000CFFECFFF800150002FFE900030015FFF7FFEC000D0010",
		INIT_51=>X"00000014FFFAFFEC000A0010FFF1FFF300120008FFEBFFFC0015FFFEFFEA0007",
		INIT_52=>X"FFEDFFFA00130000FFEB00040013FFF6FFEF000D000DFFEFFFF600130004FFEB",
		INIT_53=>X"000EFFF1FFF400110006FFEDFFFE0013FFFDFFED00070011FFF3FFF1000F000A",
		INIT_54=>X"00050011FFF6FFF1000D000BFFEFFFF800120003FFEC00010012FFF9FFEE000A",
		INIT_55=>X"FFEEFFFF0012FFFCFFEE0008000FFFF3FFF3000F0008FFEEFFFB0012FFFFFFED",
		INIT_56=>X"000AFFF0FFF900110001FFEE00020011FFF9FFF0000A000CFFF1FFF600100005",
		INIT_57=>X"0008000DFFF3FFF5000E0007FFEFFFFD0011FFFEFFEE0005000FFFF6FFF2000D",
		INIT_58=>X"FFEF00030010FFF8FFF1000B000BFFF1FFF700100004FFEE00000011FFFBFFF0",
		INIT_59=>X"0005FFEFFFFE0010FFFDFFEF0006000EFFF5FFF3000D0008FFF0FFFA00100000",
		INIT_5A=>X"000B000AFFF1FFF9000F0002FFEF00010010FFFAFFF10009000CFFF3FFF6000E",
		INIT_5B=>X"FFF00007000DFFF5FFF4000D0007FFF0FFFC0010FFFFFFEF0004000FFFF7FFF2",
		INIT_5C=>X"0001FFEF0002000FFFF9FFF10009000BFFF3FFF7000E0004FFEFFFFF0010FFFC",
		INIT_5D=>X"000D0006FFF0FFFD0010FFFEFFF00005000EFFF7FFF3000B0009FFF1FFFA000F",
		INIT_5E=>X"FFF2000A000AFFF3FFF8000E0003FFF00000000FFFFBFFF10007000CFFF4FFF5",
		INIT_5F=>X"FFFDFFF00005000EFFF6FFF4000C0008FFF1FFFB000F0000FFF00003000FFFF9",
		INIT_60=>X"000F0003FFF00000000FFFFBFFF10008000CFFF4FFF6000E0005FFF0FFFD0010",
		INIT_61=>X"FFF4000C0007FFF1FFFB000F0000FFF00003000EFFF8FFF3000A000AFFF2FFF9",
		INIT_62=>X"FFFAFFF10009000BFFF3FFF7000E0005FFF0FFFE0010FFFDFFF00006000DFFF5",
		INIT_63=>X"0010FFFFFFEF0004000EFFF7FFF3000B0009FFF1FFF9000F0002FFEF0001000F",
		INIT_64=>X"FFF7000F0004FFEFFFFF0010FFFCFFF00007000DFFF4FFF5000D0007FFF0FFFC",
		INIT_65=>X"FFF6FFF3000C0009FFF1FFFA00100001FFEF0002000FFFF9FFF1000A000BFFF2",
		INIT_66=>X"0010FFFAFFF00008000DFFF3FFF5000E0006FFEFFFFD0010FFFEFFEF0005000E",
		INIT_67=>X"FFFB00110000FFEE00040010FFF7FFF1000B000BFFF1FFF800100003FFEF0000",
		INIT_68=>X"FFF2FFF6000F0005FFEEFFFE0011FFFDFFEF0007000EFFF5FFF3000D0008FFF0",
		INIT_69=>X"0010FFF6FFF1000C000AFFF0FFF900110002FFEE00010011FFF9FFF0000A000D",
		INIT_6A=>X"FFFF0012FFFBFFEE0008000FFFF3FFF3000F0008FFEEFFFC0012FFFFFFEE0005",
		INIT_6B=>X"FFEEFFF900120001FFEC00030012FFF8FFEF000B000DFFF1FFF600110005FFED",
		INIT_6C=>X"000FFFF1FFF300110007FFEDFFFD0013FFFEFFED00060011FFF4FFF1000E000A",
		INIT_6D=>X"00040013FFF6FFEF000D000DFFEFFFF600130004FFEB00000013FFFAFFED000A",
		INIT_6E=>X"FFEAFFFE0015FFFCFFEB00080012FFF3FFF10010000AFFECFFFA00140000FFEB",
		INIT_6F=>X"000DFFECFFF700150003FFE900020015FFF8FFEC000C0010FFEFFFF300130007",
		INIT_70=>X"000A0013FFF0FFF00013000AFFEAFFFA0017FFFFFFE900060014FFF4FFEE0010",
		INIT_71=>X"FFE600030017FFF6FFEA000F0011FFECFFF300160006FFE8FFFF0017FFFAFFE9",
		INIT_72=>X"000AFFE6FFFB001AFFFDFFE600080017FFF1FFEC0013000EFFE9FFF700180002",
		INIT_73=>X"00120013FFE8FFF2001A0006FFE40000001BFFF8FFE6000D0015FFECFFEF0017",
		INIT_74=>X"FFE2000B001AFFEDFFEA0017000FFFE4FFF7001D0001FFE20006001BFFF3FFE8",
		INIT_75=>X"0005FFDE00020020FFF5FFE200120018FFE8FFED001C000BFFE1FFFC001FFFFB",
		INIT_76=>X"001E0011FFDDFFF70024FFFFFFDC00090020FFEEFFE400180015FFE2FFF20020",
		INIT_77=>X"FFDB0018001DFFE0FFEA0024000BFFD9FFFE0026FFF8FFDB0010001FFFE7FFE6",
		INIT_78=>X"FFFCFFD2000E0029FFE7FFDD00210019FFD9FFF0002A0004FFD500050028FFF0",
		INIT_79=>X"0032000CFFCA00000033FFF2FFD000190028FFDDFFE000290014FFD1FFF7002F",
		INIT_7A=>X"FFD100310021FFC6FFED003C0003FFC4000B0037FFE6FFCF00240026FFD2FFE6",
		INIT_7B=>X"FFE6FFB8002A003BFFC8FFD40041001AFFBAFFF70046FFF6FFBD0019003AFFD8",
		INIT_7C=>X"006AFFFFFF9A0019005BFFD0FFB30040003AFFB3FFDA0053000FFFAB00050050",
		INIT_7D=>X"FFAB008B002DFF71FFF70089FFE6FF8300360068FFB1FFAF005E0036FF98FFE5",
		INIT_7E=>X"FF5BFF2100C80098FF25FFA900DB001AFF2F001900BBFFBAFF620066007AFF81",
		INIT_7F=>X"1435FD76F9AF0274034BFDACFE25022600F6FE0FFFA701B1FFE6FE92006C0126",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_13,
		DOPADOP=>dopadop_13,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_14: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"0C3C3C3CF0F0F0C3C3C30F0F0F3C3C3C30F0F0F3C3C3CF0F0F0C3C3C3CF0F0F0",
		INITP_01=>X"F0F3C3C3CF0F0F0C3C3C3CF0F0F0C3C3C30F0F0F3C3C3C30F0F0F3C3C3CF0F0F",
		INITP_02=>X"0F0F3C3C3C30F0F0F3C3C3CF0F0F0C3C3C3CF0F0F0C3C3C30F0F0F3C3C3C30F0",
		INITP_03=>X"F0F0F0C3C3C30F0F0F3C3C3C30F0F0F3C3C3CF0F0F0C3C3C3CF0F0F0C3C3C30F",
		INITP_04=>X"C30F0F0C3C3C3CF0F0F0C3C3C3CF0F0F3C3C3C30F0F0F3C3C3C30F0F0C3C3C3C",
		INITP_05=>X"3C30F0F0F3C3C3C30F0F0C3C3C3CF0F0F0C3C3C3CF0F0F3C3C3C30F0F0F3C3C3",
		INITP_06=>X"C3C3CF0F0F3C3C3C30F0F0F3C3C3C30F0F0C3C3C3CF0F0F0C3C3C3CF0F0F3C3C",
		INITP_07=>X"3C3C3CF0F0F0C3C3C3CF0F0F3C3C3C30F0F0F3C3C3C30F0F0C3C3C3CF0F0F0C3",
		INITP_08=>X"33CC33CC330CF30CF30CF30CF30CC33CC33CC33CC33CC330CF30CF30CF30CF30",
		INITP_09=>X"0CF30CF30CF30CF30CC33CC33CC33CC33CC330CF30CF30CF30CF30CC33CC33CC",
		INITP_0A=>X"F30CF30CF33CC33CC33CC33CC330CF30CF30CF30CF30CC33CC33CC33CC33CC33",
		INITP_0B=>X"3CC33CC33CC33CC33CCF30CF30CF30CF30CF33CC33CC33CC33CC33CCF30CF30C",
		INITP_0C=>X"C33CC33CCF30CF30CF30CF30CF33CC33CC33CC33CC33CCF30CF30CF30CF30CF3",
		INITP_0D=>X"30CF30CF30CF30CF30CC33CC33CC33CC33CC330CF30CF30CF30CF33CC33CC33C",
		INITP_0E=>X"CF30CF30CC33CC33CC33CC33CC330CF30CF30CF30CF30CC33CC33CC33CC33CC3",
		INITP_0F=>X"33CC33CC33CC33CC330CF30CF30CF30CF30CC33CC33CC33CC33CC330CF30CF30",
		INIT_00=>X"006CFE92FFE601B1FFA7FE0F00F60226FE25FDAC034B0274F9AFFD7614352290",
		INIT_01=>X"007A0066FF62FFBA00BB0019FF2F001A00DBFFA9FF25009800C8FF21FF5B0126",
		INIT_02=>X"FF980036005EFFAFFFB100680036FF83FFE60089FFF7FF71002D008BFFABFF81",
		INIT_03=>X"0005FFAB000F0053FFDAFFB3003A0040FFB3FFD0005B0019FF9AFFFF006AFFE5",
		INIT_04=>X"003A0019FFBDFFF60046FFF7FFBA001A0041FFD4FFC8003B002AFFB8FFE60050",
		INIT_05=>X"FFD200260024FFCFFFE60037000BFFC40003003CFFEDFFC600210031FFD1FFD8",
		INIT_06=>X"FFF7FFD100140029FFE0FFDD00280019FFD0FFF200330000FFCA000C0032FFE6",
		INIT_07=>X"00280005FFD50004002AFFF0FFD900190021FFDDFFE70029000EFFD2FFFC002F",
		INIT_08=>X"FFE7001F0010FFDBFFF80026FFFEFFD9000B0024FFEAFFE0001D0018FFDBFFF0",
		INIT_09=>X"FFF2FFE200150018FFE4FFEE00200009FFDCFFFF0024FFF7FFDD0011001EFFE6",
		INIT_0A=>X"001FFFFCFFE1000B001CFFEDFFE800180012FFE2FFF500200002FFDE00050020",
		INIT_0B=>X"FFF3001B0006FFE20001001DFFF7FFE4000F0017FFEAFFED001A000BFFE2FFFB",
		INIT_0C=>X"FFEFFFEC0015000DFFE6FFF8001B0000FFE40006001AFFF2FFE800130012FFE8",
		INIT_0D=>X"0018FFF7FFE9000E0013FFECFFF100170008FFE6FFFD001AFFFBFFE6000A0017",
		INIT_0E=>X"FFFA0017FFFFFFE800060016FFF3FFEC0011000FFFEAFFF600170003FFE60002",
		INIT_0F=>X"FFEEFFF400140006FFE9FFFF0017FFFAFFEA000A0013FFF0FFF00013000AFFE9",
		INIT_10=>X"0013FFF3FFEF0010000CFFECFFF800150002FFE900030015FFF7FFEC000D0010",
		INIT_11=>X"00000014FFFAFFEC000A0010FFF1FFF300120008FFEBFFFC0015FFFEFFEA0007",
		INIT_12=>X"FFEDFFFA00130000FFEB00040013FFF6FFEF000D000DFFEFFFF600130004FFEB",
		INIT_13=>X"000EFFF1FFF400110006FFEDFFFE0013FFFDFFED00070011FFF3FFF1000F000A",
		INIT_14=>X"00050011FFF6FFF1000D000BFFEFFFF800120003FFEC00010012FFF9FFEE000A",
		INIT_15=>X"FFEEFFFF0012FFFCFFEE0008000FFFF3FFF3000F0008FFEEFFFB0012FFFFFFED",
		INIT_16=>X"000AFFF0FFF900110001FFEE00020011FFF9FFF0000A000CFFF1FFF600100005",
		INIT_17=>X"0008000DFFF3FFF5000E0007FFEFFFFD0011FFFEFFEE0005000FFFF6FFF2000D",
		INIT_18=>X"FFEF00030010FFF8FFF1000B000BFFF1FFF700100004FFEE00000011FFFBFFF0",
		INIT_19=>X"0005FFEFFFFE0010FFFDFFEF0006000EFFF5FFF3000D0008FFF0FFFA00100000",
		INIT_1A=>X"000B000AFFF1FFF9000F0002FFEF00010010FFFAFFF10009000CFFF3FFF6000E",
		INIT_1B=>X"FFF00007000DFFF5FFF4000D0007FFF0FFFC0010FFFFFFEF0004000FFFF7FFF2",
		INIT_1C=>X"0001FFEF0002000FFFF9FFF10009000BFFF3FFF7000E0004FFEFFFFF0010FFFC",
		INIT_1D=>X"000D0006FFF0FFFD0010FFFEFFF00005000EFFF7FFF3000B0009FFF1FFFA000F",
		INIT_1E=>X"FFF2000A000AFFF3FFF8000E0003FFF00000000FFFFBFFF10007000CFFF4FFF5",
		INIT_1F=>X"FFFDFFF00005000EFFF6FFF4000C0008FFF1FFFB000F0000FFF00003000FFFF9",
		INIT_20=>X"000F0003FFF00000000FFFFBFFF10008000CFFF4FFF6000E0005FFF0FFFD0010",
		INIT_21=>X"FFF4000C0007FFF1FFFB000F0000FFF00003000EFFF8FFF3000A000AFFF2FFF9",
		INIT_22=>X"FFFAFFF10009000BFFF3FFF7000E0005FFF0FFFE0010FFFDFFF00006000DFFF5",
		INIT_23=>X"0010FFFFFFEF0004000EFFF7FFF3000B0009FFF1FFF9000F0002FFEF0001000F",
		INIT_24=>X"FFF7000F0004FFEFFFFF0010FFFCFFF00007000DFFF4FFF5000D0007FFF0FFFC",
		INIT_25=>X"FFF6FFF3000C0009FFF1FFFA00100001FFEF0002000FFFF9FFF1000A000BFFF2",
		INIT_26=>X"0010FFFAFFF00008000DFFF3FFF5000E0006FFEFFFFD0010FFFEFFEF0005000E",
		INIT_27=>X"FFFB00110000FFEE00040010FFF7FFF1000B000BFFF1FFF800100003FFEF0000",
		INIT_28=>X"FFF2FFF6000F0005FFEEFFFE0011FFFDFFEF0007000EFFF5FFF3000D0008FFF0",
		INIT_29=>X"0010FFF6FFF1000C000AFFF0FFF900110002FFEE00010011FFF9FFF0000A000D",
		INIT_2A=>X"FFFF0012FFFBFFEE0008000FFFF3FFF3000F0008FFEEFFFC0012FFFFFFEE0005",
		INIT_2B=>X"FFEEFFF900120001FFEC00030012FFF8FFEF000B000DFFF1FFF600110005FFED",
		INIT_2C=>X"000FFFF1FFF300110007FFEDFFFD0013FFFEFFED00060011FFF4FFF1000E000A",
		INIT_2D=>X"00040013FFF6FFEF000D000DFFEFFFF600130004FFEB00000013FFFAFFED000A",
		INIT_2E=>X"FFEAFFFE0015FFFCFFEB00080012FFF3FFF10010000AFFECFFFA00140000FFEB",
		INIT_2F=>X"000DFFECFFF700150003FFE900020015FFF8FFEC000C0010FFEFFFF300130007",
		INIT_30=>X"000A0013FFF0FFF00013000AFFEAFFFA0017FFFFFFE900060014FFF4FFEE0010",
		INIT_31=>X"FFE600030017FFF6FFEA000F0011FFECFFF300160006FFE8FFFF0017FFFAFFE9",
		INIT_32=>X"000AFFE6FFFB001AFFFDFFE600080017FFF1FFEC0013000EFFE9FFF700180002",
		INIT_33=>X"00120013FFE8FFF2001A0006FFE40000001BFFF8FFE6000D0015FFECFFEF0017",
		INIT_34=>X"FFE2000B001AFFEDFFEA0017000FFFE4FFF7001D0001FFE20006001BFFF3FFE8",
		INIT_35=>X"0005FFDE00020020FFF5FFE200120018FFE8FFED001C000BFFE1FFFC001FFFFB",
		INIT_36=>X"001E0011FFDDFFF70024FFFFFFDC00090020FFEEFFE400180015FFE2FFF20020",
		INIT_37=>X"FFDB0018001DFFE0FFEA0024000BFFD9FFFE0026FFF8FFDB0010001FFFE7FFE6",
		INIT_38=>X"FFFCFFD2000E0029FFE7FFDD00210019FFD9FFF0002A0004FFD500050028FFF0",
		INIT_39=>X"0032000CFFCA00000033FFF2FFD000190028FFDDFFE000290014FFD1FFF7002F",
		INIT_3A=>X"FFD100310021FFC6FFED003C0003FFC4000B0037FFE6FFCF00240026FFD2FFE6",
		INIT_3B=>X"FFE6FFB8002A003BFFC8FFD40041001AFFBAFFF70046FFF6FFBD0019003AFFD8",
		INIT_3C=>X"006AFFFFFF9A0019005BFFD0FFB30040003AFFB3FFDA0053000FFFAB00050050",
		INIT_3D=>X"FFAB008B002DFF71FFF70089FFE6FF8300360068FFB1FFAF005E0036FF98FFE5",
		INIT_3E=>X"FF5BFF2100C80098FF25FFA900DB001AFF2F001900BBFFBAFF620066007AFF81",
		INIT_3F=>X"1435FD76F9AF0274034BFDACFE25022600F6FE0FFFA701B1FFE6FE92006C0126",
		INIT_40=>X"FEC80163FF3DFF910194FE020143006FFDA8035EFD71FF900519F5D20E173070",
		INIT_41=>X"FF58008BFFE2FF9600BDFF550033006BFF2600D3FFAEFF9300FFFEF3007D006D",
		INIT_42=>X"FF93003E0014FF9F0078FFB2FFF30062FF7A005E0001FF9A0095FF8D000C0067",
		INIT_43=>X"FFB90014002BFFAC004EFFE3FFD80057FFA800260022FFA50061FFCEFFE3005D",
		INIT_44=>X"FFD7FFF80034FFBA002F0001FFCD0049FFC900050030FFB3003EFFF3FFD10050",
		INIT_45=>X"FFEEFFE70035FFCB00160014FFCA0038FFE3FFEF0035FFC20022000CFFCA0041",
		INIT_46=>X"0001FFDD0030FFDB00020020FFCD0028FFF8FFE10033FFD3000C001BFFCB0030",
		INIT_47=>X"000FFFD90028FFECFFF30025FFD500170008FFDA002CFFE4FFFA0023FFD1001F",
		INIT_48=>X"0018FFDA001DFFFAFFE90026FFDF00080014FFD90023FFF3FFED0026FFDA0010",
		INIT_49=>X"001DFFDE00120007FFE30022FFEAFFFB001BFFDC00180001FFE50024FFE40001",
		INIT_4A=>X"001EFFE500060010FFE1001CFFF6FFF1001EFFE2000C000CFFE1001FFFF0FFF6",
		INIT_4B=>X"001CFFEEFFFC0016FFE200130001FFEA001EFFEA00010014FFE10017FFFCFFED",
		INIT_4C=>X"0017FFF8FFF30019FFE7000A000AFFE6001AFFF3FFF70018FFE4000E0006FFE8",
		INIT_4D=>X"00100001FFED0019FFED00000011FFE60014FFFCFFF0001AFFEA0005000EFFE5",
		INIT_4E=>X"00080009FFE90016FFF5FFF80015FFE8000C0005FFEB0018FFF1FFFC0013FFE6",
		INIT_4F=>X"0000000FFFE90011FFFDFFF10016FFED0004000CFFE90014FFF9FFF40016FFEA",
		INIT_50=>X"FFF90013FFEB000A0005FFED0015FFF3FFFC0011FFE9000E0001FFEF0016FFF0",
		INIT_51=>X"FFF30014FFEF0003000BFFEB0012FFFAFFF50014FFEC00070008FFEC0014FFF6",
		INIT_52=>X"FFEF0013FFF4FFFC0010FFEB000C0001FFF00014FFF10000000EFFEB000FFFFD",
		INIT_53=>X"FFED0010FFFBFFF60012FFEE00060007FFED0012FFF7FFF90011FFEC00090004",
		INIT_54=>X"FFED000B0001FFF10012FFF20000000DFFED000EFFFEFFF40012FFF00003000A",
		INIT_55=>X"FFEF00060007FFEF0010FFF8FFF90010FFEE00080004FFF00012FFF5FFFC000E",
		INIT_56=>X"FFF3FFFF000CFFEE000DFFFEFFF40011FFF10002000AFFEE000FFFFBFFF70011",
		INIT_57=>X"FFF9FFFA000FFFEF00080004FFF10011FFF6FFFC000EFFEE000A0001FFF20011",
		INIT_58=>X"FFFEFFF50010FFF200020009FFEF000EFFFBFFF70010FFF000050007FFEF0010",
		INIT_59=>X"0004FFF10010FFF6FFFC000DFFEF000A0001FFF30010FFF4FFFF000BFFEF000C",
		INIT_5A=>X"0009FFEF000DFFFCFFF7000FFFF100050007FFF0000FFFF9FFFA000FFFF00007",
		INIT_5B=>X"000DFFEF00090001FFF30010FFF4FFFF000BFFEF000CFFFEFFF50010FFF20002",
		INIT_5C=>X"000FFFF100040007FFF0000EFFF9FFFA000EFFF000070004FFF1000FFFF7FFFC",
		INIT_5D=>X"0010FFF5FFFF000BFFEF000BFFFFFFF50010FFF300020009FFF0000DFFFCFFF7",
		INIT_5E=>X"000EFFF9FFFA000EFFF000070004FFF2000FFFF7FFFC000DFFF000090001FFF3",
		INIT_5F=>X"000BFFFFFFF5000FFFF300020009FFF0000DFFFCFFF7000FFFF100040007FFF0",
		INIT_60=>X"00070004FFF1000FFFF7FFFC000DFFF000090002FFF3000FFFF5FFFF000BFFF0",
		INIT_61=>X"00010009FFF0000DFFFCFFF7000FFFF200040007FFF0000EFFFAFFF9000EFFF0",
		INIT_62=>X"FFFC000DFFF000090002FFF30010FFF5FFFF000BFFEF000BFFFFFFF50010FFF3",
		INIT_63=>X"FFF7000FFFF100040007FFF0000EFFFAFFF9000EFFF000070004FFF1000FFFF7",
		INIT_64=>X"FFF20010FFF5FFFE000CFFEF000BFFFFFFF40010FFF300010009FFEF000DFFFC",
		INIT_65=>X"FFF0000FFFFAFFF9000FFFF000070005FFF1000FFFF7FFFC000DFFEF00090002",
		INIT_66=>X"FFEF000BFFFFFFF40010FFF30001000AFFEF000DFFFCFFF60010FFF100040007",
		INIT_67=>X"FFEF00070005FFF00010FFF7FFFB000EFFEF00090002FFF20010FFF5FFFE000C",
		INIT_68=>X"FFF20001000AFFEE000EFFFCFFF60011FFF100040008FFEF000FFFFAFFF90010",
		INIT_69=>X"FFF7FFFB000FFFEE000A0002FFF10011FFF4FFFE000DFFEE000CFFFFFFF30011",
		INIT_6A=>X"FFFCFFF50012FFF000040008FFEE0010FFF9FFF80010FFEF00070006FFEF0011",
		INIT_6B=>X"0003FFF00012FFF4FFFE000EFFED000D0000FFF20012FFF10001000BFFED000E",
		INIT_6C=>X"0009FFEC0011FFF9FFF70012FFED00070006FFEE0012FFF6FFFB0010FFED000A",
		INIT_6D=>X"000FFFEB000E0000FFF10014FFF00001000CFFEB0010FFFCFFF40013FFEF0004",
		INIT_6E=>X"0014FFEC00080007FFEC0014FFF5FFFA0012FFEB000B0003FFEF0014FFF3FFFD",
		INIT_6F=>X"0016FFEF0001000EFFE90011FFFCFFF30015FFED0005000AFFEB0013FFF9FFF6",
		INIT_70=>X"0016FFF4FFF90014FFE9000C0004FFED0016FFF1FFFD0011FFE9000F0000FFF0",
		INIT_71=>X"0013FFFCFFF10018FFEB0005000CFFE80015FFF8FFF50016FFE900090008FFEA",
		INIT_72=>X"000E0005FFEA001AFFF0FFFC0014FFE600110000FFED0019FFED00010010FFE6",
		INIT_73=>X"0006000EFFE40018FFF7FFF3001AFFE6000A000AFFE70019FFF3FFF80017FFE5",
		INIT_74=>X"FFFC0017FFE100140001FFEA001EFFEA00010013FFE20016FFFCFFEE001CFFE8",
		INIT_75=>X"FFF0001FFFE1000C000CFFE2001EFFF1FFF6001CFFE100100006FFE5001EFFED",
		INIT_76=>X"FFE40024FFE500010018FFDC001BFFFBFFEA0022FFE300070012FFDE001DFFF6",
		INIT_77=>X"FFDA0026FFEDFFF30023FFD900140008FFDF0026FFE9FFFA001DFFDA00180001",
		INIT_78=>X"FFD10023FFFAFFE4002CFFDA00080017FFD50025FFF3FFEC0028FFD9000F0010",
		INIT_79=>X"FFCB001B000CFFD30033FFE1FFF80028FFCD00200002FFDB0030FFDD0001001F",
		INIT_7A=>X"FFCA000C0022FFC20035FFEFFFE30038FFCA00140016FFCB0035FFE7FFEE0030",
		INIT_7B=>X"FFD1FFF3003EFFB300300005FFC90049FFCD0001002FFFBA0034FFF8FFD70041",
		INIT_7C=>X"FFE3FFCE0061FFA500220026FFA80057FFD8FFE3004EFFAC002B0014FFB90050",
		INIT_7D=>X"000CFF8D0095FF9A0001005EFF7A0062FFF3FFB20078FF9F0014003EFF93005D",
		INIT_7E=>X"007DFEF300FFFF93FFAE00D3FF26006B0033FF5500BDFF96FFE2008BFF580067",
		INIT_7F=>X"0E17F5D20519FF90FD71035EFDA8006F0143FE020194FF91FF3D0163FEC8006D",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_14,
		DOPADOP=>dopadop_14,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_15: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"33CC33CC330CF30CF30CF30CF30CC33CC33CC33CC33CC330CF30CF30CF30CF30",
		INITP_01=>X"0CF30CF30CF30CF30CC33CC33CC33CC33CC330CF30CF30CF30CF30CC33CC33CC",
		INITP_02=>X"F30CF30CF33CC33CC33CC33CC330CF30CF30CF30CF30CC33CC33CC33CC33CC33",
		INITP_03=>X"3CC33CC33CC33CC33CCF30CF30CF30CF30CF33CC33CC33CC33CC33CCF30CF30C",
		INITP_04=>X"C33CC33CCF30CF30CF30CF30CF33CC33CC33CC33CC33CCF30CF30CF30CF30CF3",
		INITP_05=>X"30CF30CF30CF30CF30CC33CC33CC33CC33CC330CF30CF30CF30CF33CC33CC33C",
		INITP_06=>X"CF30CF30CC33CC33CC33CC33CC330CF30CF30CF30CF30CC33CC33CC33CC33CC3",
		INITP_07=>X"33CC33CC33CC33CC330CF30CF30CF30CF30CC33CC33CC33CC33CC330CF30CF30",
		INITP_08=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC",
		INITP_09=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0A=>X"000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0B=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_0C=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_0D=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0F=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_00=>X"FEC80163FF3DFF910194FE020143006FFDA8035EFD71FF900519F5D20E173070",
		INIT_01=>X"FF58008BFFE2FF9600BDFF550033006BFF2600D3FFAEFF9300FFFEF3007D006D",
		INIT_02=>X"FF93003E0014FF9F0078FFB2FFF30062FF7A005E0001FF9A0095FF8D000C0067",
		INIT_03=>X"FFB90014002BFFAC004EFFE3FFD80057FFA800260022FFA50061FFCEFFE3005D",
		INIT_04=>X"FFD7FFF80034FFBA002F0001FFCD0049FFC900050030FFB3003EFFF3FFD10050",
		INIT_05=>X"FFEEFFE70035FFCB00160014FFCA0038FFE3FFEF0035FFC20022000CFFCA0041",
		INIT_06=>X"0001FFDD0030FFDB00020020FFCD0028FFF8FFE10033FFD3000C001BFFCB0030",
		INIT_07=>X"000FFFD90028FFECFFF30025FFD500170008FFDA002CFFE4FFFA0023FFD1001F",
		INIT_08=>X"0018FFDA001DFFFAFFE90026FFDF00080014FFD90023FFF3FFED0026FFDA0010",
		INIT_09=>X"001DFFDE00120007FFE30022FFEAFFFB001BFFDC00180001FFE50024FFE40001",
		INIT_0A=>X"001EFFE500060010FFE1001CFFF6FFF1001EFFE2000C000CFFE1001FFFF0FFF6",
		INIT_0B=>X"001CFFEEFFFC0016FFE200130001FFEA001EFFEA00010014FFE10017FFFCFFED",
		INIT_0C=>X"0017FFF8FFF30019FFE7000A000AFFE6001AFFF3FFF70018FFE4000E0006FFE8",
		INIT_0D=>X"00100001FFED0019FFED00000011FFE60014FFFCFFF0001AFFEA0005000EFFE5",
		INIT_0E=>X"00080009FFE90016FFF5FFF80015FFE8000C0005FFEB0018FFF1FFFC0013FFE6",
		INIT_0F=>X"0000000FFFE90011FFFDFFF10016FFED0004000CFFE90014FFF9FFF40016FFEA",
		INIT_10=>X"FFF90013FFEB000A0005FFED0015FFF3FFFC0011FFE9000E0001FFEF0016FFF0",
		INIT_11=>X"FFF30014FFEF0003000BFFEB0012FFFAFFF50014FFEC00070008FFEC0014FFF6",
		INIT_12=>X"FFEF0013FFF4FFFC0010FFEB000C0001FFF00014FFF10000000EFFEB000FFFFD",
		INIT_13=>X"FFED0010FFFBFFF60012FFEE00060007FFED0012FFF7FFF90011FFEC00090004",
		INIT_14=>X"FFED000B0001FFF10012FFF20000000DFFED000EFFFEFFF40012FFF00003000A",
		INIT_15=>X"FFEF00060007FFEF0010FFF8FFF90010FFEE00080004FFF00012FFF5FFFC000E",
		INIT_16=>X"FFF3FFFF000CFFEE000DFFFEFFF40011FFF10002000AFFEE000FFFFBFFF70011",
		INIT_17=>X"FFF9FFFA000FFFEF00080004FFF10011FFF6FFFC000EFFEE000A0001FFF20011",
		INIT_18=>X"FFFEFFF50010FFF200020009FFEF000EFFFBFFF70010FFF000050007FFEF0010",
		INIT_19=>X"0004FFF10010FFF6FFFC000DFFEF000A0001FFF30010FFF4FFFF000BFFEF000C",
		INIT_1A=>X"0009FFEF000DFFFCFFF7000FFFF100050007FFF0000FFFF9FFFA000FFFF00007",
		INIT_1B=>X"000DFFEF00090001FFF30010FFF4FFFF000BFFEF000CFFFEFFF50010FFF20002",
		INIT_1C=>X"000FFFF100040007FFF0000EFFF9FFFA000EFFF000070004FFF1000FFFF7FFFC",
		INIT_1D=>X"0010FFF5FFFF000BFFEF000BFFFFFFF50010FFF300020009FFF0000DFFFCFFF7",
		INIT_1E=>X"000EFFF9FFFA000EFFF000070004FFF2000FFFF7FFFC000DFFF000090001FFF3",
		INIT_1F=>X"000BFFFFFFF5000FFFF300020009FFF0000DFFFCFFF7000FFFF100040007FFF0",
		INIT_20=>X"00070004FFF1000FFFF7FFFC000DFFF000090002FFF3000FFFF5FFFF000BFFF0",
		INIT_21=>X"00010009FFF0000DFFFCFFF7000FFFF200040007FFF0000EFFFAFFF9000EFFF0",
		INIT_22=>X"FFFC000DFFF000090002FFF30010FFF5FFFF000BFFEF000BFFFFFFF50010FFF3",
		INIT_23=>X"FFF7000FFFF100040007FFF0000EFFFAFFF9000EFFF000070004FFF1000FFFF7",
		INIT_24=>X"FFF20010FFF5FFFE000CFFEF000BFFFFFFF40010FFF300010009FFEF000DFFFC",
		INIT_25=>X"FFF0000FFFFAFFF9000FFFF000070005FFF1000FFFF7FFFC000DFFEF00090002",
		INIT_26=>X"FFEF000BFFFFFFF40010FFF30001000AFFEF000DFFFCFFF60010FFF100040007",
		INIT_27=>X"FFEF00070005FFF00010FFF7FFFB000EFFEF00090002FFF20010FFF5FFFE000C",
		INIT_28=>X"FFF20001000AFFEE000EFFFCFFF60011FFF100040008FFEF000FFFFAFFF90010",
		INIT_29=>X"FFF7FFFB000FFFEE000A0002FFF10011FFF4FFFE000DFFEE000CFFFFFFF30011",
		INIT_2A=>X"FFFCFFF50012FFF000040008FFEE0010FFF9FFF80010FFEF00070006FFEF0011",
		INIT_2B=>X"0003FFF00012FFF4FFFE000EFFED000D0000FFF20012FFF10001000BFFED000E",
		INIT_2C=>X"0009FFEC0011FFF9FFF70012FFED00070006FFEE0012FFF6FFFB0010FFED000A",
		INIT_2D=>X"000FFFEB000E0000FFF10014FFF00001000CFFEB0010FFFCFFF40013FFEF0004",
		INIT_2E=>X"0014FFEC00080007FFEC0014FFF5FFFA0012FFEB000B0003FFEF0014FFF3FFFD",
		INIT_2F=>X"0016FFEF0001000EFFE90011FFFCFFF30015FFED0005000AFFEB0013FFF9FFF6",
		INIT_30=>X"0016FFF4FFF90014FFE9000C0004FFED0016FFF1FFFD0011FFE9000F0000FFF0",
		INIT_31=>X"0013FFFCFFF10018FFEB0005000CFFE80015FFF8FFF50016FFE900090008FFEA",
		INIT_32=>X"000E0005FFEA001AFFF0FFFC0014FFE600110000FFED0019FFED00010010FFE6",
		INIT_33=>X"0006000EFFE40018FFF7FFF3001AFFE6000A000AFFE70019FFF3FFF80017FFE5",
		INIT_34=>X"FFFC0017FFE100140001FFEA001EFFEA00010013FFE20016FFFCFFEE001CFFE8",
		INIT_35=>X"FFF0001FFFE1000C000CFFE2001EFFF1FFF6001CFFE100100006FFE5001EFFED",
		INIT_36=>X"FFE40024FFE500010018FFDC001BFFFBFFEA0022FFE300070012FFDE001DFFF6",
		INIT_37=>X"FFDA0026FFEDFFF30023FFD900140008FFDF0026FFE9FFFA001DFFDA00180001",
		INIT_38=>X"FFD10023FFFAFFE4002CFFDA00080017FFD50025FFF3FFEC0028FFD9000F0010",
		INIT_39=>X"FFCB001B000CFFD30033FFE1FFF80028FFCD00200002FFDB0030FFDD0001001F",
		INIT_3A=>X"FFCA000C0022FFC20035FFEFFFE30038FFCA00140016FFCB0035FFE7FFEE0030",
		INIT_3B=>X"FFD1FFF3003EFFB300300005FFC90049FFCD0001002FFFBA0034FFF8FFD70041",
		INIT_3C=>X"FFE3FFCE0061FFA500220026FFA80057FFD8FFE3004EFFAC002B0014FFB90050",
		INIT_3D=>X"000CFF8D0095FF9A0001005EFF7A0062FFF3FFB20078FF9F0014003EFF93005D",
		INIT_3E=>X"007DFEF300FFFF93FFAE00D3FF26006B0033FF5500BDFF96FFE2008BFF580067",
		INIT_3F=>X"0E17F5D20519FF90FD71035EFDA8006F0143FE020194FF91FF3D0163FEC8006D",
		INIT_40=>X"FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD03FD0",
		INIT_41=>X"FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0",
		INIT_42=>X"FFD1FFD1FFD1FFD1FFD1FFD1FFD1FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0",
		INIT_43=>X"FFD2FFD2FFD2FFD2FFD2FFD2FFD1FFD1FFD1FFD1FFD1FFD1FFD1FFD1FFD1FFD1",
		INIT_44=>X"FFD3FFD3FFD3FFD3FFD3FFD3FFD3FFD3FFD2FFD2FFD2FFD2FFD2FFD2FFD2FFD2",
		INIT_45=>X"FFD5FFD5FFD5FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD3FFD3FFD3",
		INIT_46=>X"FFD7FFD7FFD6FFD6FFD6FFD6FFD6FFD6FFD6FFD6FFD5FFD5FFD5FFD5FFD5FFD5",
		INIT_47=>X"FFD9FFD9FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD7FFD7FFD7FFD7FFD7FFD7",
		INIT_48=>X"FFDBFFDBFFDBFFDBFFDAFFDAFFDAFFDAFFDAFFDAFFDAFFD9FFD9FFD9FFD9FFD9",
		INIT_49=>X"FFDEFFDDFFDDFFDDFFDDFFDDFFDDFFDCFFDCFFDCFFDCFFDCFFDCFFDCFFDBFFDB",
		INIT_4A=>X"FFE0FFE0FFE0FFE0FFE0FFDFFFDFFFDFFFDFFFDFFFDFFFDEFFDEFFDEFFDEFFDE",
		INIT_4B=>X"FFE3FFE3FFE3FFE3FFE2FFE2FFE2FFE2FFE2FFE1FFE1FFE1FFE1FFE1FFE1FFE0",
		INIT_4C=>X"FFE6FFE6FFE6FFE5FFE5FFE5FFE5FFE5FFE5FFE4FFE4FFE4FFE4FFE4FFE3FFE3",
		INIT_4D=>X"FFE9FFE9FFE9FFE8FFE8FFE8FFE8FFE8FFE8FFE7FFE7FFE7FFE7FFE7FFE6FFE6",
		INIT_4E=>X"FFECFFECFFECFFECFFEBFFEBFFEBFFEBFFEBFFEAFFEAFFEAFFEAFFEAFFE9FFE9",
		INIT_4F=>X"FFEFFFEFFFEFFFEFFFEFFFEEFFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEC",
		INIT_50=>X"FFF2FFF2FFF2FFF2FFF2FFF1FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFF0FFF0",
		INIT_51=>X"FFF6FFF5FFF5FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3FFF3FFF3FFF3",
		INIT_52=>X"FFF9FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6",
		INIT_53=>X"FFFCFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9",
		INIT_54=>X"FFFEFFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFC",
		INIT_55=>X"0001000100010001000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_56=>X"0004000300030003000300030003000300020002000200020002000200010001",
		INIT_57=>X"0006000600060006000500050005000500050005000500040004000400040004",
		INIT_58=>X"0008000800080008000800070007000700070007000700070007000600060006",
		INIT_59=>X"000A000A000A000A000A00090009000900090009000900090009000800080008",
		INIT_5A=>X"000C000C000B000B000B000B000B000B000B000B000B000B000A000A000A000A",
		INIT_5B=>X"000D000D000D000D000D000D000D000C000C000C000C000C000C000C000C000C",
		INIT_5C=>X"000E000E000E000E000E000E000E000E000E000D000D000D000D000D000D000D",
		INIT_5D=>X"000F000F000F000F000F000F000F000F000E000E000E000E000E000E000E000E",
		INIT_5E=>X"000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F",
		INIT_5F=>X"000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F",
		INIT_60=>X"000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F0010",
		INIT_61=>X"000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F000F",
		INIT_62=>X"000E000E000E000E000E000E000E000F000F000F000F000F000F000F000F000F",
		INIT_63=>X"000D000D000D000D000D000D000E000E000E000E000E000E000E000E000E000E",
		INIT_64=>X"000C000C000C000C000C000C000C000C000D000D000D000D000D000D000D000D",
		INIT_65=>X"000A000A000A000B000B000B000B000B000B000B000B000B000B000C000C000C",
		INIT_66=>X"0008000800090009000900090009000900090009000A000A000A000A000A000A",
		INIT_67=>X"0006000600070007000700070007000700070007000800080008000800080008",
		INIT_68=>X"0004000400040004000500050005000500050005000500060006000600060006",
		INIT_69=>X"0001000200020002000200020002000300030003000300030003000300040004",
		INIT_6A=>X"FFFFFFFFFFFFFFFFFFFF00000000000000000000000000010001000100010001",
		INIT_6B=>X"FFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFEFFFEFFFF",
		INIT_6C=>X"FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFCFFFC",
		INIT_6D=>X"FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF9FFF9",
		INIT_6E=>X"FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF5FFF6FFF6",
		INIT_6F=>X"FFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2FFF2FFF3",
		INIT_70=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEFFFEFFFF0",
		INIT_71=>X"FFE9FFEAFFEAFFEAFFEAFFEAFFEBFFEBFFEBFFEBFFEBFFECFFECFFECFFECFFEC",
		INIT_72=>X"FFE6FFE7FFE7FFE7FFE7FFE7FFE8FFE8FFE8FFE8FFE8FFE8FFE9FFE9FFE9FFE9",
		INIT_73=>X"FFE3FFE4FFE4FFE4FFE4FFE4FFE5FFE5FFE5FFE5FFE5FFE5FFE6FFE6FFE6FFE6",
		INIT_74=>X"FFE1FFE1FFE1FFE1FFE1FFE1FFE2FFE2FFE2FFE2FFE2FFE3FFE3FFE3FFE3FFE3",
		INIT_75=>X"FFDEFFDEFFDEFFDEFFDFFFDFFFDFFFDFFFDFFFDFFFE0FFE0FFE0FFE0FFE0FFE0",
		INIT_76=>X"FFDBFFDCFFDCFFDCFFDCFFDCFFDCFFDCFFDDFFDDFFDDFFDDFFDDFFDDFFDEFFDE",
		INIT_77=>X"FFD9FFD9FFD9FFD9FFDAFFDAFFDAFFDAFFDAFFDAFFDAFFDBFFDBFFDBFFDBFFDB",
		INIT_78=>X"FFD7FFD7FFD7FFD7FFD7FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD8FFD9FFD9FFD9",
		INIT_79=>X"FFD5FFD5FFD5FFD5FFD5FFD6FFD6FFD6FFD6FFD6FFD6FFD6FFD6FFD7FFD7FFD7",
		INIT_7A=>X"FFD3FFD3FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD4FFD5FFD5FFD5FFD5",
		INIT_7B=>X"FFD2FFD2FFD2FFD2FFD2FFD2FFD2FFD3FFD3FFD3FFD3FFD3FFD3FFD3FFD3FFD3",
		INIT_7C=>X"FFD1FFD1FFD1FFD1FFD1FFD1FFD1FFD1FFD1FFD2FFD2FFD2FFD2FFD2FFD2FFD2",
		INIT_7D=>X"FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD1FFD1FFD1FFD1FFD1FFD1FFD1FFD1",
		INIT_7E=>X"FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0",
		INIT_7F=>X"FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0FFD0",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_15,
		DOPADOP=>dopadop_15,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
end arch;
