library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity filter_table is
	port(
		clk:  in  std_logic;
		addr: in  std_logic_vector(14 downto 0);
		data: out signed(17 downto 0)
	);
end filter_table;

architecture arch of filter_table is
	signal addr_d:  std_logic_vector(14 downto 11);
	signal addrardaddr:   std_logic_vector(15 downto 0);
	signal doado_00:  std_logic_vector(31 downto 0);
	signal dopadop_00: std_logic_vector(3 downto 0);
	signal doado_01:  std_logic_vector(31 downto 0);
	signal dopadop_01: std_logic_vector(3 downto 0);
	signal doado_02:  std_logic_vector(31 downto 0);
	signal dopadop_02: std_logic_vector(3 downto 0);
	signal doado_03:  std_logic_vector(31 downto 0);
	signal dopadop_03: std_logic_vector(3 downto 0);
	signal doado_04:  std_logic_vector(31 downto 0);
	signal dopadop_04: std_logic_vector(3 downto 0);
	signal doado_05:  std_logic_vector(31 downto 0);
	signal dopadop_05: std_logic_vector(3 downto 0);
	signal doado_06:  std_logic_vector(31 downto 0);
	signal dopadop_06: std_logic_vector(3 downto 0);
	signal doado_07:  std_logic_vector(31 downto 0);
	signal dopadop_07: std_logic_vector(3 downto 0);
	signal doado_08:  std_logic_vector(31 downto 0);
	signal dopadop_08: std_logic_vector(3 downto 0);
	signal doado_09:  std_logic_vector(31 downto 0);
	signal dopadop_09: std_logic_vector(3 downto 0);
	signal doado_10:  std_logic_vector(31 downto 0);
	signal dopadop_10: std_logic_vector(3 downto 0);
	signal doado_11:  std_logic_vector(31 downto 0);
	signal dopadop_11: std_logic_vector(3 downto 0);
	signal doado_12:  std_logic_vector(31 downto 0);
	signal dopadop_12: std_logic_vector(3 downto 0);
	signal doado_13:  std_logic_vector(31 downto 0);
	signal dopadop_13: std_logic_vector(3 downto 0);
	signal doado_14:  std_logic_vector(31 downto 0);
	signal dopadop_14: std_logic_vector(3 downto 0);
	signal doado_15:  std_logic_vector(31 downto 0);
	signal dopadop_15: std_logic_vector(3 downto 0);
begin
	addrardaddr(15)<='1';
	addrardaddr(14 downto 4)<=addr(10 downto 0);
	addrardaddr(3 downto 0)<=b"0000";
	process(clk)
	begin
		if (rising_edge(clk)) then
			addr_d<=addr(14 downto 11);
		end if;
	end process;
	with addr_d select data(15 downto 0)<=
		signed(doado_00(15 downto 0)) when b"0000",
		signed(doado_01(15 downto 0)) when b"0001",
		signed(doado_02(15 downto 0)) when b"0010",
		signed(doado_03(15 downto 0)) when b"0011",
		signed(doado_04(15 downto 0)) when b"0100",
		signed(doado_05(15 downto 0)) when b"0101",
		signed(doado_06(15 downto 0)) when b"0110",
		signed(doado_07(15 downto 0)) when b"0111",
		signed(doado_08(15 downto 0)) when b"1000",
		signed(doado_09(15 downto 0)) when b"1001",
		signed(doado_10(15 downto 0)) when b"1010",
		signed(doado_11(15 downto 0)) when b"1011",
		signed(doado_12(15 downto 0)) when b"1100",
		signed(doado_13(15 downto 0)) when b"1101",
		signed(doado_14(15 downto 0)) when b"1110",
		signed(doado_15(15 downto 0)) when others;
	with addr_d select data(17 downto 16)<=
		signed(dopadop_00(1 downto 0)) when b"0000",
		signed(dopadop_01(1 downto 0)) when b"0001",
		signed(dopadop_02(1 downto 0)) when b"0010",
		signed(dopadop_03(1 downto 0)) when b"0011",
		signed(dopadop_04(1 downto 0)) when b"0100",
		signed(dopadop_05(1 downto 0)) when b"0101",
		signed(dopadop_06(1 downto 0)) when b"0110",
		signed(dopadop_07(1 downto 0)) when b"0111",
		signed(dopadop_08(1 downto 0)) when b"1000",
		signed(dopadop_09(1 downto 0)) when b"1001",
		signed(dopadop_10(1 downto 0)) when b"1010",
		signed(dopadop_11(1 downto 0)) when b"1011",
		signed(dopadop_12(1 downto 0)) when b"1100",
		signed(dopadop_13(1 downto 0)) when b"1101",
		signed(dopadop_14(1 downto 0)) when b"1110",
		signed(dopadop_15(1 downto 0)) when others;
	mem_00: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_01=>X"0000000000000000000000000000000000000000000000000000000FFFFFFFFF",
		INITP_02=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000",
		INITP_04=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_05=>X"0000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_06=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_08=>X"000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_09=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_0A=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000",
		INITP_0B=>X"000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0C=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_0D=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000",
		INITP_0E=>X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0F=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_00=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_01=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_02=>X"FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_03=>X"FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_04=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9",
		INIT_05=>X"FFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFA",
		INIT_06=>X"FFFDFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFB",
		INIT_07=>X"FFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFD",
		INIT_08=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFE",
		INIT_09=>X"00010001000100000000000000000000000000000000000000000000FFFFFFFF",
		INIT_0A=>X"0002000200020002000200020002000100010001000100010001000100010001",
		INIT_0B=>X"0003000300030003000300030003000300030003000300030002000200020002",
		INIT_0C=>X"0005000500050004000400040004000400040004000400040004000400040004",
		INIT_0D=>X"0006000600060006000600050005000500050005000500050005000500050005",
		INIT_0E=>X"0007000700070007000700060006000600060006000600060006000600060006",
		INIT_0F=>X"0008000700070007000700070007000700070007000700070007000700070007",
		INIT_10=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_11=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_12=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_13=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_14=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_15=>X"0007000700070007000700070007000700070007000700080008000800080008",
		INIT_16=>X"0006000600060006000600060006000600070007000700070007000700070007",
		INIT_17=>X"0005000500050005000500050005000500050006000600060006000600060006",
		INIT_18=>X"0003000400040004000400040004000400040004000400040005000500050005",
		INIT_19=>X"0002000200020002000200020003000300030003000300030003000300030003",
		INIT_1A=>X"0000000000000001000100010001000100010001000100010002000200020002",
		INIT_1B=>X"FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000",
		INIT_1C=>X"FFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFE",
		INIT_1D=>X"FFFBFFFBFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFD",
		INIT_1E=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFB",
		INIT_1F=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_20=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_21=>X"FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_22=>X"FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5",
		INIT_23=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4",
		INIT_24=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3",
		INIT_25=>X"FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3",
		INIT_26=>X"FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF2FFF2",
		INIT_27=>X"FFF4FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3",
		INIT_28=>X"FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4",
		INIT_29=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5",
		INIT_2A=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF6FFF6",
		INIT_2B=>X"FFFBFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8",
		INIT_2C=>X"FFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFB",
		INIT_2D=>X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFE",
		INIT_2E=>X"0004000400030003000300030003000200020002000200010001000100010001",
		INIT_2F=>X"0007000700070007000700060006000600060005000500050005000400040004",
		INIT_30=>X"000B000B000B000B000A000A000A000A00090009000900090008000800080008",
		INIT_31=>X"000F000F000F000F000E000E000E000E000D000D000D000D000C000C000C000C",
		INIT_32=>X"0014001300130013001300120012001200120011001100110010001000100010",
		INIT_33=>X"0018001800170017001700160016001600160015001500150015001400140014",
		INIT_34=>X"001C001C001B001B001B001B001A001A001A001A001900190019001900180018",
		INIT_35=>X"002000200020001F001F001F001F001E001E001E001E001D001D001D001C001C",
		INIT_36=>X"0024002400240023002300230023002200220022002200210021002100210020",
		INIT_37=>X"0028002700270027002700270026002600260026002500250025002500240024",
		INIT_38=>X"002B002B002B002B002A002A002A002A00290029002900290029002800280028",
		INIT_39=>X"002E002E002E002E002E002D002D002D002D002D002C002C002C002C002C002B",
		INIT_3A=>X"0031003100310031003000300030003000300030002F002F002F002F002F002E",
		INIT_3B=>X"0033003300330033003300330032003200320032003200320032003100310031",
		INIT_3C=>X"0035003500350035003500350034003400340034003400340034003400340033",
		INIT_3D=>X"0036003600360036003600360036003600360036003600360035003500350035",
		INIT_3E=>X"0037003700370037003700370037003700370037003700370037003700370036",
		INIT_3F=>X"0038003700370037003700370037003700370037003700370037003700370037",
		INIT_40=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_41=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_42=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_43=>X"FFFCFFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFA",
		INIT_44=>X"FFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFC",
		INIT_45=>X"000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFE",
		INIT_46=>X"0002000200020002000200010001000100010001000100010000000000000000",
		INIT_47=>X"0004000400040004000400030003000300030003000300030003000200020002",
		INIT_48=>X"0006000600060005000500050005000500050005000500050004000400040004",
		INIT_49=>X"0007000700070007000700070007000600060006000600060006000600060006",
		INIT_4A=>X"0008000800080008000800080007000700070007000700070007000700070007",
		INIT_4B=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_4C=>X"0007000700070007000800080008000800080008000800080008000800080008",
		INIT_4D=>X"0006000600060007000700070007000700070007000700070007000700070007",
		INIT_4E=>X"0005000500050005000500050005000600060006000600060006000600060006",
		INIT_4F=>X"0003000300030003000300030004000400040004000400040004000400050005",
		INIT_50=>X"0001000100010001000100010001000200020002000200020002000200030003",
		INIT_51=>X"FFFEFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000",
		INIT_52=>X"FFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFE",
		INIT_53=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFCFFFC",
		INIT_54=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFFAFFFA",
		INIT_55=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_56=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_57=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_58=>X"FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_59=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_5A=>X"FFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_5B=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFA",
		INIT_5C=>X"FFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFD",
		INIT_5D=>X"000200020002000200010001000100010001000000000000000000000000FFFF",
		INIT_5E=>X"0005000500050004000400040004000400040003000300030003000300020002",
		INIT_5F=>X"0008000700070007000700070007000600060006000600060006000500050005",
		INIT_60=>X"000A000900090009000900090009000900090008000800080008000800080008",
		INIT_61=>X"000B000B000B000B000B000B000B000B000A000A000A000A000A000A000A000A",
		INIT_62=>X"000C000C000C000C000C000C000C000C000C000B000B000B000B000B000B000B",
		INIT_63=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C",
		INIT_64=>X"000A000B000B000B000B000B000B000B000B000B000B000B000B000B000B000C",
		INIT_65=>X"00090009000900090009000900090009000A000A000A000A000A000A000A000A",
		INIT_66=>X"0006000600060006000700070007000700070007000800080008000800080008",
		INIT_67=>X"0002000300030003000300030004000400040004000500050005000500050006",
		INIT_68=>X"FFFEFFFFFFFFFFFFFFFF00000000000000000001000100010001000200020002",
		INIT_69=>X"FFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFEFFFEFFFE",
		INIT_6A=>X"FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFA",
		INIT_6B=>X"FFF2FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6",
		INIT_6C=>X"FFEFFFEFFFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2",
		INIT_6D=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEF",
		INIT_6E=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFED",
		INIT_6F=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_70=>X"FFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFECFFECFFECFFEC",
		INIT_71=>X"FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEEFFEEFFEE",
		INIT_72=>X"FFF6FFF6FFF6FFF5FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF2FFF2FFF2FFF2",
		INIT_73=>X"FFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF7FFF7FFF7",
		INIT_74=>X"00050004000400030003000200020001000100000000FFFFFFFFFFFEFFFEFFFD",
		INIT_75=>X"000E000D000C000C000B000B000A000A00090008000800070007000600060005",
		INIT_76=>X"0017001700160015001500140014001300120012001100110010000F000F000E",
		INIT_77=>X"0022002100200020001F001E001E001D001C001C001B001B001A001900190018",
		INIT_78=>X"002C002B002B002A002900290028002700270026002500250024002400230022",
		INIT_79=>X"00360035003500340034003300320032003100300030002F002E002E002D002D",
		INIT_7A=>X"003F003F003E003E003D003C003C003B003B003A003A00390038003800370037",
		INIT_7B=>X"0047004700470046004600450045004400440043004200420041004100400040",
		INIT_7C=>X"004E004E004E004D004D004C004C004B004B004B004A004A0049004900480048",
		INIT_7D=>X"0053005300530053005200520052005100510051005000500050004F004F004F",
		INIT_7E=>X"0056005600560056005600560056005500550055005500550054005400540054",
		INIT_7F=>X"0058005700570057005700570057005700570057005700570057005700570057",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_00,
		DOPADOP=>dopadop_00,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_01: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_01=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000",
		INITP_03=>X"000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_04=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000",
		INITP_06=>X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_08=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000",
		INITP_09=>X"00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0A=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000",
		INITP_0B=>X"0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFF",
		INITP_0C=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000",
		INITP_0D=>X"00000000000000000000000000000000000000000000000000000FFFFFFFFFFF",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000",
		INITP_0F=>X"0000000000000000000000000000000000000000000000000000000000003FFF",
		INIT_00=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_01=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_02=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_03=>X"FFFCFFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFA",
		INIT_04=>X"FFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFC",
		INIT_05=>X"000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFE",
		INIT_06=>X"0002000200020002000200010001000100010001000100010000000000000000",
		INIT_07=>X"0004000400040004000400030003000300030003000300030003000200020002",
		INIT_08=>X"0006000600060005000500050005000500050005000500050004000400040004",
		INIT_09=>X"0007000700070007000700070007000600060006000600060006000600060006",
		INIT_0A=>X"0008000800080008000800080007000700070007000700070007000700070007",
		INIT_0B=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_0C=>X"0007000700070007000800080008000800080008000800080008000800080008",
		INIT_0D=>X"0006000600060007000700070007000700070007000700070007000700070007",
		INIT_0E=>X"0005000500050005000500050005000600060006000600060006000600060006",
		INIT_0F=>X"0003000300030003000300030004000400040004000400040004000400050005",
		INIT_10=>X"0001000100010001000100010001000200020002000200020002000200030003",
		INIT_11=>X"FFFEFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000",
		INIT_12=>X"FFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFE",
		INIT_13=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFCFFFC",
		INIT_14=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFFAFFFA",
		INIT_15=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_16=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_17=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_18=>X"FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_19=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_1A=>X"FFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_1B=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFA",
		INIT_1C=>X"FFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFD",
		INIT_1D=>X"000200020002000200010001000100010001000000000000000000000000FFFF",
		INIT_1E=>X"0005000500050004000400040004000400040003000300030003000300020002",
		INIT_1F=>X"0008000700070007000700070007000600060006000600060006000500050005",
		INIT_20=>X"000A000900090009000900090009000900090008000800080008000800080008",
		INIT_21=>X"000B000B000B000B000B000B000B000B000A000A000A000A000A000A000A000A",
		INIT_22=>X"000C000C000C000C000C000C000C000C000C000B000B000B000B000B000B000B",
		INIT_23=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C",
		INIT_24=>X"000A000B000B000B000B000B000B000B000B000B000B000B000B000B000B000C",
		INIT_25=>X"00090009000900090009000900090009000A000A000A000A000A000A000A000A",
		INIT_26=>X"0006000600060006000700070007000700070007000800080008000800080008",
		INIT_27=>X"0002000300030003000300030004000400040004000500050005000500050006",
		INIT_28=>X"FFFEFFFFFFFFFFFFFFFF00000000000000000001000100010001000200020002",
		INIT_29=>X"FFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFEFFFEFFFE",
		INIT_2A=>X"FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFA",
		INIT_2B=>X"FFF2FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6",
		INIT_2C=>X"FFEFFFEFFFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2",
		INIT_2D=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEF",
		INIT_2E=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFED",
		INIT_2F=>X"FFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFECFFEC",
		INIT_30=>X"FFEEFFEEFFEEFFEEFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFEDFFECFFECFFECFFEC",
		INIT_31=>X"FFF1FFF1FFF1FFF1FFF0FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEEFFEEFFEE",
		INIT_32=>X"FFF6FFF6FFF6FFF5FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF3FFF2FFF2FFF2FFF2",
		INIT_33=>X"FFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF7FFF7FFF7",
		INIT_34=>X"00050004000400030003000200020001000100000000FFFFFFFFFFFEFFFEFFFD",
		INIT_35=>X"000E000D000C000C000B000B000A000A00090008000800070007000600060005",
		INIT_36=>X"0017001700160015001500140014001300120012001100110010000F000F000E",
		INIT_37=>X"0022002100200020001F001E001E001D001C001C001B001B001A001900190018",
		INIT_38=>X"002C002B002B002A002900290028002700270026002500250024002400230022",
		INIT_39=>X"00360035003500340034003300320032003100300030002F002E002E002D002D",
		INIT_3A=>X"003F003F003E003E003D003C003C003B003B003A003A00390038003800370037",
		INIT_3B=>X"0047004700470046004600450045004400440043004200420041004100400040",
		INIT_3C=>X"004E004E004E004D004D004C004C004B004B004B004A004A0049004900480048",
		INIT_3D=>X"0053005300530053005200520052005100510051005000500050004F004F004F",
		INIT_3E=>X"0056005600560056005600560056005500550055005500550054005400540054",
		INIT_3F=>X"0058005700570057005700570057005700570057005700570057005700570057",
		INIT_40=>X"0007000700070007000700070007000700070007000700070007000700070007",
		INIT_41=>X"0005000500050005000500060006000600060006000600060006000700070007",
		INIT_42=>X"0002000200020003000300030003000300040004000400040004000400050005",
		INIT_43=>X"FFFFFFFFFFFFFFFF000000000000000000000001000100010001000100020002",
		INIT_44=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFF",
		INIT_45=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFB",
		INIT_46=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9",
		INIT_47=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8",
		INIT_48=>X"FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_49=>X"FFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9",
		INIT_4A=>X"FFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFB",
		INIT_4B=>X"000200020002000100010001000100000000000000000000FFFFFFFFFFFFFFFF",
		INIT_4C=>X"0005000500050004000400040004000400040003000300030003000300020002",
		INIT_4D=>X"0007000700070007000700070006000600060006000600060006000500050005",
		INIT_4E=>X"0008000800080008000800080008000800080008000800080008000700070007",
		INIT_4F=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_50=>X"0006000600060006000600060006000700070007000700070007000700070007",
		INIT_51=>X"0002000300030003000300040004000400040004000400050005000500050005",
		INIT_52=>X"FFFFFFFFFFFF0000000000000000000000010001000100010002000200020002",
		INIT_53=>X"FFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFF",
		INIT_54=>X"FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFB",
		INIT_55=>X"FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_56=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_57=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_58=>X"FFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_59=>X"FFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFA",
		INIT_5A=>X"00020002000200010001000100010000000000000000FFFFFFFFFFFFFFFFFFFE",
		INIT_5B=>X"0006000600060005000500050005000400040004000400030003000300030002",
		INIT_5C=>X"0009000900090009000800080008000800080007000700070007000700060006",
		INIT_5D=>X"000A000A000A000A000A000A000A000A000A000A000A000A0009000900090009",
		INIT_5E=>X"000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A",
		INIT_5F=>X"0008000800080008000800080009000900090009000900090009000A000A000A",
		INIT_60=>X"0004000400040004000500050005000600060006000600060007000700070007",
		INIT_61=>X"FFFFFFFF00000000000000000001000100010002000200020003000300030003",
		INIT_62=>X"FFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFEFFFF",
		INIT_63=>X"FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFA",
		INIT_64=>X"FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF5FFF6",
		INIT_65=>X"FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3",
		INIT_66=>X"FFF4FFF4FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF2",
		INIT_67=>X"FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF4FFF4FFF4",
		INIT_68=>X"FFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_69=>X"0003000300020002000200010001000000000000FFFFFFFFFFFEFFFEFFFEFFFD",
		INIT_6A=>X"0009000900090008000800080007000700060006000600050005000400040004",
		INIT_6B=>X"000E000E000E000E000D000D000D000D000C000C000C000B000B000B000A000A",
		INIT_6C=>X"001100110011001100110011001100100010001000100010000F000F000F000F",
		INIT_6D=>X"0011001100110011001100110012001200120012001200120012001100110011",
		INIT_6E=>X"000E000E000E000F000F000F000F001000100010001000100011001100110011",
		INIT_6F=>X"00080008000800090009000A000A000B000B000B000C000C000C000D000D000D",
		INIT_70=>X"FFFF000000000001000100020002000300030004000500050006000600070007",
		INIT_71=>X"FFF5FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFBFFFCFFFDFFFDFFFEFFFE",
		INIT_72=>X"FFECFFEDFFEDFFEEFFEEFFEFFFEFFFF0FFF1FFF1FFF2FFF2FFF3FFF4FFF4FFF5",
		INIT_73=>X"FFE5FFE5FFE6FFE6FFE7FFE7FFE7FFE8FFE8FFE9FFE9FFEAFFEAFFEBFFEBFFEC",
		INIT_74=>X"FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE3FFE3FFE3FFE3FFE4FFE4FFE4FFE4FFE5",
		INIT_75=>X"FFE3FFE3FFE3FFE3FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2",
		INIT_76=>X"FFEAFFEAFFE9FFE9FFE8FFE8FFE7FFE7FFE6FFE6FFE5FFE5FFE5FFE4FFE4FFE4",
		INIT_77=>X"FFF7FFF7FFF6FFF5FFF4FFF3FFF2FFF1FFF0FFEFFFEFFFEEFFEDFFECFFECFFEB",
		INIT_78=>X"000A00080007000600050004000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF8",
		INIT_79=>X"0020001F001D001C001A0019001700160014001300120010000F000E000C000B",
		INIT_7A=>X"003800370035003400320031002F002E002C002B002900270026002400230021",
		INIT_7B=>X"0051004F004E004C004B0049004800460045004300420040003F003D003B003A",
		INIT_7C=>X"006700650064006300620060005F005E005C005B005900580057005500540052",
		INIT_7D=>X"007800770076007500740073007200710070006F006E006D006C006A00690068",
		INIT_7E=>X"00840083008300820081008100800080007F007E007D007D007C007B007A0079",
		INIT_7F=>X"0088008700870087008700870087008700870086008600860085008500850084",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_01,
		DOPADOP=>dopadop_01,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_02: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000",
		INITP_01=>X"00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_02=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000",
		INITP_03=>X"0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFF",
		INITP_04=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000",
		INITP_05=>X"00000000000000000000000000000000000000000000000000000FFFFFFFFFFF",
		INITP_06=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000",
		INITP_07=>X"0000000000000000000000000000000000000000000000000000000000003FFF",
		INITP_08=>X"000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF",
		INITP_09=>X"00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00",
		INITP_0A=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000",
		INITP_0B=>X"FFFFFFFFFFFC00000000000000000000000000000000000000000000FFFFFFFF",
		INITP_0C=>X"0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0D=>X"000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000",
		INITP_0F=>X"000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
		INIT_00=>X"0007000700070007000700070007000700070007000700070007000700070007",
		INIT_01=>X"0005000500050005000500060006000600060006000600060006000700070007",
		INIT_02=>X"0002000200020003000300030003000300040004000400040004000400050005",
		INIT_03=>X"FFFFFFFFFFFFFFFF000000000000000000000001000100010001000100020002",
		INIT_04=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFF",
		INIT_05=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFB",
		INIT_06=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9",
		INIT_07=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8",
		INIT_08=>X"FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_09=>X"FFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9",
		INIT_0A=>X"FFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFB",
		INIT_0B=>X"000200020002000100010001000100000000000000000000FFFFFFFFFFFFFFFF",
		INIT_0C=>X"0005000500050004000400040004000400040003000300030003000300020002",
		INIT_0D=>X"0007000700070007000700070006000600060006000600060006000500050005",
		INIT_0E=>X"0008000800080008000800080008000800080008000800080008000700070007",
		INIT_0F=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_10=>X"0006000600060006000600060006000700070007000700070007000700070007",
		INIT_11=>X"0002000300030003000300040004000400040004000400050005000500050005",
		INIT_12=>X"FFFFFFFFFFFF0000000000000000000000010001000100010002000200020002",
		INIT_13=>X"FFFBFFFBFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFF",
		INIT_14=>X"FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFBFFFBFFFB",
		INIT_15=>X"FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_16=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_17=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_18=>X"FFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_19=>X"FFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFA",
		INIT_1A=>X"00020002000200010001000100010000000000000000FFFFFFFFFFFFFFFFFFFE",
		INIT_1B=>X"0006000600060005000500050005000400040004000400030003000300030002",
		INIT_1C=>X"0009000900090009000800080008000800080007000700070007000700060006",
		INIT_1D=>X"000A000A000A000A000A000A000A000A000A000A000A000A0009000900090009",
		INIT_1E=>X"000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A000A",
		INIT_1F=>X"0008000800080008000800080009000900090009000900090009000A000A000A",
		INIT_20=>X"0004000400040004000500050005000600060006000600060007000700070007",
		INIT_21=>X"FFFFFFFF00000000000000000001000100010002000200020003000300030003",
		INIT_22=>X"FFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFEFFFF",
		INIT_23=>X"FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFA",
		INIT_24=>X"FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF5FFF6",
		INIT_25=>X"FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3",
		INIT_26=>X"FFF4FFF4FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF2FFF2FFF2FFF2FFF2",
		INIT_27=>X"FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF4FFF4FFF4",
		INIT_28=>X"FFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_29=>X"0003000300020002000200010001000000000000FFFFFFFFFFFEFFFEFFFEFFFD",
		INIT_2A=>X"0009000900090008000800080007000700060006000600050005000400040004",
		INIT_2B=>X"000E000E000E000E000D000D000D000D000C000C000C000B000B000B000A000A",
		INIT_2C=>X"001100110011001100110011001100100010001000100010000F000F000F000F",
		INIT_2D=>X"0011001100110011001100110012001200120012001200120012001100110011",
		INIT_2E=>X"000E000E000E000F000F000F000F001000100010001000100011001100110011",
		INIT_2F=>X"00080008000800090009000A000A000B000B000B000C000C000C000D000D000D",
		INIT_30=>X"FFFF000000000001000100020002000300030004000500050006000600070007",
		INIT_31=>X"FFF5FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFBFFFCFFFDFFFDFFFEFFFE",
		INIT_32=>X"FFECFFEDFFEDFFEEFFEEFFEFFFEFFFF0FFF1FFF1FFF2FFF2FFF3FFF4FFF4FFF5",
		INIT_33=>X"FFE5FFE5FFE6FFE6FFE7FFE7FFE7FFE8FFE8FFE9FFE9FFEAFFEAFFEBFFEBFFEC",
		INIT_34=>X"FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE3FFE3FFE3FFE3FFE4FFE4FFE4FFE4FFE5",
		INIT_35=>X"FFE3FFE3FFE3FFE3FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2FFE2",
		INIT_36=>X"FFEAFFEAFFE9FFE9FFE8FFE8FFE7FFE7FFE6FFE6FFE5FFE5FFE5FFE4FFE4FFE4",
		INIT_37=>X"FFF7FFF7FFF6FFF5FFF4FFF3FFF2FFF1FFF0FFEFFFEFFFEEFFEDFFECFFECFFEB",
		INIT_38=>X"000A00080007000600050004000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF8",
		INIT_39=>X"0020001F001D001C001A0019001700160014001300120010000F000E000C000B",
		INIT_3A=>X"003800370035003400320031002F002E002C002B002900270026002400230021",
		INIT_3B=>X"0051004F004E004C004B0049004800460045004300420040003F003D003B003A",
		INIT_3C=>X"006700650064006300620060005F005E005C005B005900580057005500540052",
		INIT_3D=>X"007800770076007500740073007200710070006F006E006D006C006A00690068",
		INIT_3E=>X"00840083008300820081008100800080007F007E007D007D007C007B007A0079",
		INIT_3F=>X"0088008700870087008700870087008700870086008600860085008500850084",
		INIT_40=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_41=>X"FFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9",
		INIT_42=>X"0000000000000000FFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFC",
		INIT_43=>X"0005000400040004000400030003000300030002000200020002000100010001",
		INIT_44=>X"0007000700070007000700070006000600060006000600060005000500050005",
		INIT_45=>X"0007000700070008000800080008000800080008000800070007000700070007",
		INIT_46=>X"0005000500050006000600060006000600070007000700070007000700070007",
		INIT_47=>X"0001000100020002000200020003000300030003000400040004000400050005",
		INIT_48=>X"FFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFFFFFFFFFFFFFF00000000000000010001",
		INIT_49=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFCFFFCFFFC",
		INIT_4A=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9",
		INIT_4B=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_4C=>X"FFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8",
		INIT_4D=>X"00000000FFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFCFFFC",
		INIT_4E=>X"0004000400040004000300030003000300020002000200010001000100010000",
		INIT_4F=>X"0008000700070007000700070007000600060006000600060005000500050005",
		INIT_50=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_51=>X"0006000600060007000700070007000700070008000800080008000800080008",
		INIT_52=>X"0002000200020003000300030004000400040004000500050005000500060006",
		INIT_53=>X"FFFDFFFDFFFDFFFEFFFEFFFEFFFFFFFFFFFF0000000000000001000100010002",
		INIT_54=>X"FFF9FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFD",
		INIT_55=>X"FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_56=>X"FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_57=>X"FFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7",
		INIT_58=>X"FFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFCFFFBFFFBFFFBFFFA",
		INIT_59=>X"0005000400040004000300030003000200020002000100010001000000000000",
		INIT_5A=>X"0009000800080008000800080007000700070007000600060006000600050005",
		INIT_5B=>X"000A000A000A000A000A000A000A000A000A0009000900090009000900090009",
		INIT_5C=>X"00080008000800080009000900090009000900090009000A000A000A000A000A",
		INIT_5D=>X"0003000300040004000500050005000500060006000600070007000700070008",
		INIT_5E=>X"FFFDFFFDFFFEFFFEFFFFFFFFFFFF000000000001000100010002000200020003",
		INIT_5F=>X"FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFCFFFD",
		INIT_60=>X"FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_61=>X"FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4",
		INIT_62=>X"FFF8FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF4",
		INIT_63=>X"FFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8",
		INIT_64=>X"00050005000400040004000300030002000200010001000000000000FFFFFFFF",
		INIT_65=>X"000B000B000A000A000A000A0009000900080008000800070007000700060006",
		INIT_66=>X"000D000D000D000D000D000D000D000D000D000D000C000C000C000C000C000B",
		INIT_67=>X"000B000C000C000C000C000D000D000D000D000D000D000D000D000D000D000D",
		INIT_68=>X"0006000600060007000700080008000900090009000A000A000A000B000B000B",
		INIT_69=>X"FFFDFFFEFFFEFFFFFFFF00000000000100020002000300030004000400050005",
		INIT_6A=>X"FFF5FFF5FFF6FFF6FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFCFFFCFFFD",
		INIT_6B=>X"FFEFFFEFFFF0FFF0FFF0FFF1FFF1FFF1FFF2FFF2FFF2FFF3FFF3FFF4FFF4FFF4",
		INIT_6C=>X"FFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEF",
		INIT_6D=>X"FFF3FFF2FFF2FFF2FFF1FFF1FFF1FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEE",
		INIT_6E=>X"FFFCFFFBFFFBFFFAFFFAFFF9FFF8FFF8FFF7FFF7FFF6FFF5FFF5FFF4FFF4FFF3",
		INIT_6F=>X"000800070006000500050004000300020002000100000000FFFFFFFEFFFDFFFD",
		INIT_70=>X"0012001100110010000F000F000E000E000D000C000C000B000A000A00090008",
		INIT_71=>X"0017001700170017001600160016001600150015001400140014001300130012",
		INIT_72=>X"0016001600160017001700170017001700170018001800180018001800170017",
		INIT_73=>X"000C000D000E000F000F00100011001100120013001300140014001500150015",
		INIT_74=>X"FFFDFFFEFFFF0000000100020003000400050006000700080009000A000B000C",
		INIT_75=>X"FFECFFEDFFEEFFEFFFF0FFF1FFF2FFF3FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFC",
		INIT_76=>X"FFDDFFDEFFDFFFE0FFE0FFE1FFE2FFE3FFE4FFE5FFE6FFE7FFE8FFE9FFEAFFEB",
		INIT_77=>X"FFD7FFD7FFD7FFD8FFD8FFD8FFD8FFD9FFD9FFD9FFDAFFDAFFDBFFDBFFDCFFDD",
		INIT_78=>X"FFDEFFDDFFDCFFDBFFDBFFDAFFDAFFD9FFD9FFD8FFD8FFD8FFD8FFD7FFD7FFD7",
		INIT_79=>X"FFF2FFF1FFEFFFEDFFECFFEAFFE9FFE7FFE6FFE5FFE4FFE3FFE1FFE0FFDFFFDE",
		INIT_7A=>X"00140012000F000D000B00080006000400020000FFFEFFFCFFFAFFF8FFF6FFF4",
		INIT_7B=>X"003F003C0039003600330031002E002B0029002600230021001E001B00190016",
		INIT_7C=>X"006B0069006600630060005E005B0058005500520050004D004A004700440041",
		INIT_7D=>X"00930091008F008C008A0088008500830080007E007B0079007600730071006E",
		INIT_7E=>X"00AE00AD00AB00AA00A900A700A600A400A200A1009F009D009B009900970095",
		INIT_7F=>X"00B800B700B700B700B700B700B600B600B500B400B400B300B200B100B000AF",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_02,
		DOPADOP=>dopadop_02,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_03: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF",
		INITP_01=>X"00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00",
		INITP_02=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000",
		INITP_03=>X"FFFFFFFFFFFC00000000000000000000000000000000000000000000FFFFFFFF",
		INITP_04=>X"0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_05=>X"000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000",
		INITP_06=>X"FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000",
		INITP_07=>X"000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
		INITP_08=>X"000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000",
		INITP_09=>X"00000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000",
		INITP_0A=>X"0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000",
		INITP_0B=>X"000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000",
		INITP_0C=>X"00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000",
		INITP_0D=>X"0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000",
		INITP_0E=>X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000",
		INITP_0F=>X"00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0",
		INIT_00=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_01=>X"FFFCFFFCFFFCFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9",
		INIT_02=>X"0000000000000000FFFFFFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFDFFFC",
		INIT_03=>X"0005000400040004000400030003000300030002000200020002000100010001",
		INIT_04=>X"0007000700070007000700070006000600060006000600060005000500050005",
		INIT_05=>X"0007000700070008000800080008000800080008000800070007000700070007",
		INIT_06=>X"0005000500050006000600060006000600070007000700070007000700070007",
		INIT_07=>X"0001000100020002000200020003000300030003000400040004000400050005",
		INIT_08=>X"FFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFFFFFFFFFFFFFF00000000000000010001",
		INIT_09=>X"FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFCFFFCFFFC",
		INIT_0A=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9",
		INIT_0B=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_0C=>X"FFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8",
		INIT_0D=>X"00000000FFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFCFFFC",
		INIT_0E=>X"0004000400040004000300030003000300020002000200010001000100010000",
		INIT_0F=>X"0008000700070007000700070007000600060006000600060005000500050005",
		INIT_10=>X"0008000800080008000800080008000800080008000800080008000800080008",
		INIT_11=>X"0006000600060007000700070007000700070008000800080008000800080008",
		INIT_12=>X"0002000200020003000300030004000400040004000500050005000500060006",
		INIT_13=>X"FFFDFFFDFFFDFFFEFFFEFFFEFFFFFFFFFFFF0000000000000001000100010002",
		INIT_14=>X"FFF9FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFCFFFCFFFCFFFD",
		INIT_15=>X"FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_16=>X"FFF7FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF6",
		INIT_17=>X"FFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7",
		INIT_18=>X"FFFFFFFFFFFFFFFEFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFCFFFBFFFBFFFBFFFA",
		INIT_19=>X"0005000400040004000300030003000200020002000100010001000000000000",
		INIT_1A=>X"0009000800080008000800080007000700070007000600060006000600050005",
		INIT_1B=>X"000A000A000A000A000A000A000A000A000A0009000900090009000900090009",
		INIT_1C=>X"00080008000800080009000900090009000900090009000A000A000A000A000A",
		INIT_1D=>X"0003000300040004000500050005000500060006000600070007000700070008",
		INIT_1E=>X"FFFDFFFDFFFEFFFEFFFFFFFFFFFF000000000001000100010002000200020003",
		INIT_1F=>X"FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFCFFFD",
		INIT_20=>X"FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF6FFF7FFF7FFF7",
		INIT_21=>X"FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4",
		INIT_22=>X"FFF8FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF4",
		INIT_23=>X"FFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF8",
		INIT_24=>X"00050005000400040004000300030002000200010001000000000000FFFFFFFF",
		INIT_25=>X"000B000B000A000A000A000A0009000900080008000800070007000700060006",
		INIT_26=>X"000D000D000D000D000D000D000D000D000D000D000C000C000C000C000C000B",
		INIT_27=>X"000B000C000C000C000C000D000D000D000D000D000D000D000D000D000D000D",
		INIT_28=>X"0006000600060007000700080008000900090009000A000A000A000B000B000B",
		INIT_29=>X"FFFDFFFEFFFEFFFFFFFF00000000000100020002000300030004000400050005",
		INIT_2A=>X"FFF5FFF5FFF6FFF6FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFCFFFCFFFD",
		INIT_2B=>X"FFEFFFEFFFF0FFF0FFF0FFF1FFF1FFF1FFF2FFF2FFF2FFF3FFF3FFF4FFF4FFF4",
		INIT_2C=>X"FFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEEFFEFFFEFFFEFFFEF",
		INIT_2D=>X"FFF3FFF2FFF2FFF2FFF1FFF1FFF1FFF0FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEE",
		INIT_2E=>X"FFFCFFFBFFFBFFFAFFFAFFF9FFF8FFF8FFF7FFF7FFF6FFF5FFF5FFF4FFF4FFF3",
		INIT_2F=>X"000800070006000500050004000300020002000100000000FFFFFFFEFFFDFFFD",
		INIT_30=>X"0012001100110010000F000F000E000E000D000C000C000B000A000A00090008",
		INIT_31=>X"0017001700170017001600160016001600150015001400140014001300130012",
		INIT_32=>X"0016001600160017001700170017001700170018001800180018001800170017",
		INIT_33=>X"000C000D000E000F000F00100011001100120013001300140014001500150015",
		INIT_34=>X"FFFDFFFEFFFF0000000100020003000400050006000700080009000A000B000C",
		INIT_35=>X"FFECFFEDFFEEFFEFFFF0FFF1FFF2FFF3FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFC",
		INIT_36=>X"FFDDFFDEFFDFFFE0FFE0FFE1FFE2FFE3FFE4FFE5FFE6FFE7FFE8FFE9FFEAFFEB",
		INIT_37=>X"FFD7FFD7FFD7FFD8FFD8FFD8FFD8FFD9FFD9FFD9FFDAFFDAFFDBFFDBFFDCFFDD",
		INIT_38=>X"FFDEFFDDFFDCFFDBFFDBFFDAFFDAFFD9FFD9FFD8FFD8FFD8FFD8FFD7FFD7FFD7",
		INIT_39=>X"FFF2FFF1FFEFFFEDFFECFFEAFFE9FFE7FFE6FFE5FFE4FFE3FFE1FFE0FFDFFFDE",
		INIT_3A=>X"00140012000F000D000B00080006000400020000FFFEFFFCFFFAFFF8FFF6FFF4",
		INIT_3B=>X"003F003C0039003600330031002E002B0029002600230021001E001B00190016",
		INIT_3C=>X"006B0069006600630060005E005B0058005500520050004D004A004700440041",
		INIT_3D=>X"00930091008F008C008A0088008500830080007E007B0079007600730071006E",
		INIT_3E=>X"00AE00AD00AB00AA00A900A700A600A400A200A1009F009D009B009900970095",
		INIT_3F=>X"00B800B700B700B700B700B700B600B600B500B400B400B300B200B100B000AF",
		INIT_40=>X"0005000500060006000600060006000700070007000700070007000700070007",
		INIT_41=>X"FFFF000000000000000100010002000200020003000300030004000400040005",
		INIT_42=>X"FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFEFFFEFFFEFFFF",
		INIT_43=>X"FFF8FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9",
		INIT_44=>X"FFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_45=>X"000100000000FFFFFFFFFFFFFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFCFFFBFFFB",
		INIT_46=>X"0006000600060005000500050004000400040003000300030002000200010001",
		INIT_47=>X"0008000800080008000800080008000800070007000700070007000700070006",
		INIT_48=>X"0004000400050005000500050006000600060006000700070007000700070007",
		INIT_49=>X"FFFDFFFEFFFEFFFFFFFF00000000000000010001000200020002000300030004",
		INIT_4A=>X"FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFCFFFDFFFD",
		INIT_4B=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8",
		INIT_4C=>X"FFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8",
		INIT_4D=>X"0002000200020001000100000000FFFFFFFFFFFFFFFEFFFEFFFDFFFDFFFCFFFC",
		INIT_4E=>X"0007000700070007000600060006000600050005000500040004000400030003",
		INIT_4F=>X"0007000800080008000800080008000800080008000800080008000800080008",
		INIT_50=>X"0003000300030004000400050005000500060006000600060007000700070007",
		INIT_51=>X"FFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFFFFFF0000000000010001000100020002",
		INIT_52=>X"FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFAFFFBFFFBFFFB",
		INIT_53=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_54=>X"FFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_55=>X"00040004000300030003000200020001000100000000FFFFFFFFFFFEFFFEFFFD",
		INIT_56=>X"0009000900080008000800080008000700070007000700060006000500050005",
		INIT_57=>X"0008000800080008000800090009000900090009000900090009000900090009",
		INIT_58=>X"0001000200020003000300040004000400050005000600060006000700070007",
		INIT_59=>X"FFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFEFFFEFFFFFFFF000000000001",
		INIT_5A=>X"FFF5FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9",
		INIT_5B=>X"FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5",
		INIT_5C=>X"FFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8",
		INIT_5D=>X"000700060006000500050004000400030003000200020001000100000000FFFF",
		INIT_5E=>X"000B000A000A000A000A000A000A000A00090009000900090008000800080007",
		INIT_5F=>X"0008000800080009000900090009000A000A000A000A000A000A000B000B000B",
		INIT_60=>X"FFFF000000000001000200020003000300040004000500050006000600070007",
		INIT_61=>X"FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFEFFFF",
		INIT_62=>X"FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF6FFF6FFF6",
		INIT_63=>X"FFF8FFF7FFF7FFF6FFF6FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3FFF3",
		INIT_64=>X"000100000000FFFFFFFEFFFEFFFDFFFDFFFCFFFBFFFBFFFAFFFAFFF9FFF8FFF8",
		INIT_65=>X"000A000A00090009000800080007000700060006000500040004000300020002",
		INIT_66=>X"000D000D000D000D000D000D000D000D000D000D000C000C000C000B000B000B",
		INIT_67=>X"0008000800090009000A000A000B000B000B000C000C000C000D000D000D000D",
		INIT_68=>X"FFFCFFFDFFFEFFFEFFFF00000001000100020003000400040005000600060007",
		INIT_69=>X"FFF2FFF3FFF3FFF4FFF4FFF5FFF5FFF6FFF7FFF7FFF8FFF9FFF9FFFAFFFBFFFB",
		INIT_6A=>X"FFF0FFF0FFF0FFF0FFEFFFEFFFF0FFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF2",
		INIT_6B=>X"FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF1FFF1FFF1FFF0FFF0",
		INIT_6C=>X"0005000400030002000200010000FFFFFFFEFFFDFFFCFFFBFFFBFFFAFFF9FFF8",
		INIT_6D=>X"00100010000F000F000E000E000D000C000C000B000A00090008000800070006",
		INIT_6E=>X"0012001200120013001300130013001300130013001200120012001200110011",
		INIT_6F=>X"000800080009000A000B000C000D000D000E000F000F00100010001100110012",
		INIT_70=>X"FFF6FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF0000000100020004000500060007",
		INIT_71=>X"FFE9FFEAFFEAFFEBFFECFFECFFEDFFEEFFEFFFF0FFF0FFF1FFF2FFF3FFF4FFF5",
		INIT_72=>X"FFE9FFE8FFE8FFE8FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE8FFE8FFE8FFE9",
		INIT_73=>X"FFF7FFF6FFF5FFF4FFF3FFF2FFF0FFEFFFEEFFEEFFEDFFECFFEBFFEAFFEAFFE9",
		INIT_74=>X"000E000D000B000A0009000700060004000300010000FFFEFFFDFFFCFFFAFFF9",
		INIT_75=>X"001F001F001E001D001C001C001B001A00180017001600150014001200110010",
		INIT_76=>X"001E001F00200020002100210021002200220022002200210021002100200020",
		INIT_77=>X"00080009000B000D000F0011001200140015001700180019001B001C001D001E",
		INIT_78=>X"FFE5FFE7FFE9FFEBFFEDFFF0FFF2FFF4FFF6FFF9FFFBFFFDFFFF000100030006",
		INIT_79=>X"FFCAFFCBFFCCFFCDFFCEFFD0FFD1FFD3FFD5FFD6FFD8FFDAFFDCFFDEFFE0FFE2",
		INIT_7A=>X"FFCCFFCBFFCAFFC9FFC8FFC7FFC7FFC6FFC6FFC6FFC6FFC6FFC7FFC7FFC8FFC9",
		INIT_7B=>X"FFF8FFF4FFF0FFECFFE9FFE5FFE2FFDFFFDDFFDAFFD7FFD5FFD3FFD1FFCFFFCD",
		INIT_7C=>X"00470041003B00360030002B00260021001C00170012000D000900040000FFFC",
		INIT_7D=>X"00A2009D00970092008C00860080007B0075006F00690063005D00580052004C",
		INIT_7E=>X"00EC00E800E400E100DD00D900D400D000CB00C700C200BD00B800B200AD00A8",
		INIT_7F=>X"01080107010701060106010501030102010000FE00FC00FA00F800F500F200EF",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_03,
		DOPADOP=>dopadop_03,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_04: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000",
		INITP_01=>X"00000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000",
		INITP_02=>X"0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000",
		INITP_03=>X"000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000",
		INITP_04=>X"00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000",
		INITP_05=>X"0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000",
		INITP_06=>X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000",
		INITP_07=>X"00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0",
		INITP_08=>X"0000000000FFFFFFFFFFFFFFFFFFFFFC0000000000000000000003FFFFFFFFFF",
		INITP_09=>X"FFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFF000000000000",
		INITP_0A=>X"0000000FFFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFF",
		INITP_0B=>X"FFFFFC0000000000000000000003FFFFFFFFFFFFFFFFFFFFFC00000000000000",
		INITP_0C=>X"00003FFFFFFFFFFFFFFFFFFFFF0000000000000000000000FFFFFFFFFFFFFFFF",
		INITP_0D=>X"FFF0000000000000000000000FFFFFFFFFFFFFFFFFFFFFC00000000000000000",
		INITP_0E=>X"03FFFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFF",
		INITP_0F=>X"0000000000000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000000000",
		INIT_00=>X"0005000500060006000600060006000700070007000700070007000700070007",
		INIT_01=>X"FFFF000000000000000100010002000200020003000300030004000400040005",
		INIT_02=>X"FFF9FFFAFFFAFFFAFFFBFFFBFFFBFFFCFFFCFFFCFFFDFFFDFFFEFFFEFFFEFFFF",
		INIT_03=>X"FFF8FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9",
		INIT_04=>X"FFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_05=>X"000100000000FFFFFFFFFFFFFFFEFFFEFFFDFFFDFFFDFFFCFFFCFFFCFFFBFFFB",
		INIT_06=>X"0006000600060005000500050004000400040003000300030002000200010001",
		INIT_07=>X"0008000800080008000800080008000800070007000700070007000700070006",
		INIT_08=>X"0004000400050005000500050006000600060006000700070007000700070007",
		INIT_09=>X"FFFDFFFEFFFEFFFFFFFF00000000000000010001000200020002000300030004",
		INIT_0A=>X"FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFCFFFDFFFD",
		INIT_0B=>X"FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8",
		INIT_0C=>X"FFFCFFFBFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8",
		INIT_0D=>X"0002000200020001000100000000FFFFFFFFFFFFFFFEFFFEFFFDFFFDFFFCFFFC",
		INIT_0E=>X"0007000700070007000600060006000600050005000500040004000400030003",
		INIT_0F=>X"0007000800080008000800080008000800080008000800080008000800080008",
		INIT_10=>X"0003000300030004000400050005000500060006000600060007000700070007",
		INIT_11=>X"FFFCFFFCFFFDFFFDFFFDFFFEFFFEFFFFFFFF0000000000010001000100020002",
		INIT_12=>X"FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFAFFFBFFFBFFFB",
		INIT_13=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_14=>X"FFFDFFFDFFFCFFFCFFFBFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF9FFF8FFF8FFF8",
		INIT_15=>X"00040004000300030003000200020001000100000000FFFFFFFFFFFEFFFEFFFD",
		INIT_16=>X"0009000900080008000800080008000700070007000700060006000500050005",
		INIT_17=>X"0008000800080008000800090009000900090009000900090009000900090009",
		INIT_18=>X"0001000200020003000300040004000400050005000600060006000700070007",
		INIT_19=>X"FFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFEFFFEFFFFFFFF000000000001",
		INIT_1A=>X"FFF5FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9",
		INIT_1B=>X"FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5",
		INIT_1C=>X"FFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8",
		INIT_1D=>X"000700060006000500050004000400030003000200020001000100000000FFFF",
		INIT_1E=>X"000B000A000A000A000A000A000A000A00090009000900090008000800080007",
		INIT_1F=>X"0008000800080009000900090009000A000A000A000A000A000A000B000B000B",
		INIT_20=>X"FFFF000000000001000200020003000300040004000500050006000600070007",
		INIT_21=>X"FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFEFFFF",
		INIT_22=>X"FFF3FFF3FFF3FFF3FFF3FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF6FFF6FFF6",
		INIT_23=>X"FFF8FFF7FFF7FFF6FFF6FFF5FFF5FFF5FFF4FFF4FFF4FFF4FFF4FFF3FFF3FFF3",
		INIT_24=>X"000100000000FFFFFFFEFFFEFFFDFFFDFFFCFFFBFFFBFFFAFFFAFFF9FFF8FFF8",
		INIT_25=>X"000A000A00090009000800080007000700060006000500040004000300020002",
		INIT_26=>X"000D000D000D000D000D000D000D000D000D000D000C000C000C000B000B000B",
		INIT_27=>X"0008000800090009000A000A000B000B000B000C000C000C000D000D000D000D",
		INIT_28=>X"FFFCFFFDFFFEFFFEFFFF00000001000100020003000400040005000600060007",
		INIT_29=>X"FFF2FFF3FFF3FFF4FFF4FFF5FFF5FFF6FFF7FFF7FFF8FFF9FFF9FFFAFFFBFFFB",
		INIT_2A=>X"FFF0FFF0FFF0FFF0FFEFFFEFFFF0FFF0FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF2",
		INIT_2B=>X"FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF1FFF1FFF1FFF0FFF0",
		INIT_2C=>X"0005000400030002000200010000FFFFFFFEFFFDFFFCFFFBFFFBFFFAFFF9FFF8",
		INIT_2D=>X"00100010000F000F000E000E000D000C000C000B000A00090008000800070006",
		INIT_2E=>X"0012001200120013001300130013001300130013001200120012001200110011",
		INIT_2F=>X"000800080009000A000B000C000D000D000E000F000F00100010001100110012",
		INIT_30=>X"FFF6FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF0000000100020004000500060007",
		INIT_31=>X"FFE9FFEAFFEAFFEBFFECFFECFFEDFFEEFFEFFFF0FFF0FFF1FFF2FFF3FFF4FFF5",
		INIT_32=>X"FFE9FFE8FFE8FFE8FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE8FFE8FFE8FFE9",
		INIT_33=>X"FFF7FFF6FFF5FFF4FFF3FFF2FFF0FFEFFFEEFFEEFFEDFFECFFEBFFEAFFEAFFE9",
		INIT_34=>X"000E000D000B000A0009000700060004000300010000FFFEFFFDFFFCFFFAFFF9",
		INIT_35=>X"001F001F001E001D001C001C001B001A00180017001600150014001200110010",
		INIT_36=>X"001E001F00200020002100210021002200220022002200210021002100200020",
		INIT_37=>X"00080009000B000D000F0011001200140015001700180019001B001C001D001E",
		INIT_38=>X"FFE5FFE7FFE9FFEBFFEDFFF0FFF2FFF4FFF6FFF9FFFBFFFDFFFF000100030006",
		INIT_39=>X"FFCAFFCBFFCCFFCDFFCEFFD0FFD1FFD3FFD5FFD6FFD8FFDAFFDCFFDEFFE0FFE2",
		INIT_3A=>X"FFCCFFCBFFCAFFC9FFC8FFC7FFC7FFC6FFC6FFC6FFC6FFC6FFC7FFC7FFC8FFC9",
		INIT_3B=>X"FFF8FFF4FFF0FFECFFE9FFE5FFE2FFDFFFDDFFDAFFD7FFD5FFD3FFD1FFCFFFCD",
		INIT_3C=>X"00470041003B00360030002B00260021001C00170012000D000900040000FFFC",
		INIT_3D=>X"00A2009D00970092008C00860080007B0075006F00690063005D00580052004C",
		INIT_3E=>X"00EC00E800E400E100DD00D900D400D000CB00C700C200BD00B800B200AD00A8",
		INIT_3F=>X"01080107010701060106010501030102010000FE00FC00FA00F800F500F200EF",
		INIT_40=>X"FFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_41=>X"00050004000400030003000200020001000100000000FFFFFFFEFFFEFFFDFFFD",
		INIT_42=>X"0007000700070007000800080007000700070007000700070006000600060005",
		INIT_43=>X"0000000100010002000300030004000400050005000500060006000600070007",
		INIT_44=>X"FFF8FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFEFFFFFFFF0000",
		INIT_45=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_46=>X"0001000100000000FFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9",
		INIT_47=>X"0007000700070007000700060006000600050005000400040003000300020002",
		INIT_48=>X"0004000500050006000600060007000700070007000700080008000800080008",
		INIT_49=>X"FFFBFFFCFFFCFFFDFFFDFFFEFFFFFFFF00000000000100020002000300030004",
		INIT_4A=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFB",
		INIT_4B=>X"FFFDFFFDFFFCFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF8FFF8FFF8FFF8FFF7FFF7",
		INIT_4C=>X"000600050005000500040004000300020002000100010000FFFFFFFFFFFEFFFE",
		INIT_4D=>X"0007000700080008000800080008000800080008000800070007000700070006",
		INIT_4E=>X"FFFF000000010001000200020003000300040004000500050006000600070007",
		INIT_4F=>X"FFF8FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFEFFFF",
		INIT_50=>X"FFF9FFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_51=>X"00020002000100010000FFFFFFFFFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFA",
		INIT_52=>X"0008000800080008000800080007000700070006000600050005000400040003",
		INIT_53=>X"0004000400050005000600060007000700070008000800080008000800080008",
		INIT_54=>X"FFFAFFFAFFFBFFFCFFFCFFFDFFFDFFFEFFFFFFFF000000010001000200030003",
		INIT_55=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9",
		INIT_56=>X"FFFEFFFDFFFDFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF7",
		INIT_57=>X"00080007000700060006000500040004000300030002000100010000FFFFFFFF",
		INIT_58=>X"0008000800080009000900090009000900090009000900090009000800080008",
		INIT_59=>X"FFFEFFFFFFFF0000000100020002000300040004000500050006000600070007",
		INIT_5A=>X"FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFD",
		INIT_5B=>X"FFF9FFF8FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF6",
		INIT_5C=>X"0004000400030002000100010000FFFFFFFEFFFEFFFDFFFCFFFBFFFBFFFAFFFA",
		INIT_5D=>X"000A000A000A000A000A000A0009000900090008000800070007000600060005",
		INIT_5E=>X"000300040005000600060007000700080008000900090009000A000A000A000A",
		INIT_5F=>X"FFF8FFF8FFF9FFF9FFFAFFFBFFFCFFFCFFFDFFFEFFFF00000000000100020003",
		INIT_60=>X"FFF5FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6FFF7",
		INIT_61=>X"FFFFFFFEFFFDFFFCFFFCFFFBFFFAFFF9FFF9FFF8FFF7FFF7FFF6FFF6FFF5FFF5",
		INIT_62=>X"000A000A00090009000800080007000600060005000400030002000100010000",
		INIT_63=>X"0009000A000A000B000B000B000C000C000C000C000C000C000C000B000B000B",
		INIT_64=>X"FFFCFFFDFFFEFFFF000000010002000200030004000500060007000700080009",
		INIT_65=>X"FFF2FFF2FFF3FFF3FFF3FFF4FFF4FFF5FFF6FFF6FFF7FFF8FFF9FFF9FFFAFFFB",
		INIT_66=>X"FFF8FFF7FFF6FFF6FFF5FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2",
		INIT_67=>X"000800070006000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9",
		INIT_68=>X"000E000E000E000E000E000E000E000D000D000D000C000B000B000A00090008",
		INIT_69=>X"0003000400050006000700080009000A000B000B000C000D000D000D000E000E",
		INIT_6A=>X"FFF3FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFDFFFEFFFF000000010002",
		INIT_6B=>X"FFF1FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFF0FFF0FFF1FFF1FFF2",
		INIT_6C=>X"00010000FFFEFFFDFFFCFFFBFFF9FFF8FFF7FFF6FFF5FFF4FFF3FFF2FFF2FFF1",
		INIT_6D=>X"001100110010000F000E000E000D000C000B0009000800070006000500030002",
		INIT_6E=>X"000D000E000F0010001000110011001200120012001300130012001200120012",
		INIT_6F=>X"FFF7FFF9FFFAFFFCFFFDFFFF0000000200030005000600070009000A000B000C",
		INIT_70=>X"FFE9FFE9FFEAFFEAFFEBFFEBFFECFFEDFFEEFFEFFFF0FFF1FFF2FFF3FFF5FFF6",
		INIT_71=>X"FFF5FFF4FFF2FFF1FFF0FFEFFFEEFFEDFFECFFEBFFEBFFEAFFEAFFE9FFE9FFE9",
		INIT_72=>X"0010000F000D000B000A00080006000500030001FFFFFFFEFFFCFFFAFFF8FFF7",
		INIT_73=>X"001A001A001A001B001B001A001A001A00190018001700160015001400130012",
		INIT_74=>X"0003000500070009000B000D000F001000120013001500160017001800190019",
		INIT_75=>X"FFE3FFE5FFE6FFE8FFEAFFECFFEEFFF0FFF2FFF4FFF6FFF8FFFAFFFDFFFF0001",
		INIT_76=>X"FFE2FFE0FFDFFFDFFFDEFFDDFFDDFFDDFFDDFFDDFFDEFFDEFFDFFFE0FFE1FFE2",
		INIT_77=>X"000800050002FFFFFFFCFFF9FFF6FFF4FFF1FFEFFFECFFEAFFE8FFE6FFE5FFE3",
		INIT_78=>X"002D002C002A00290027002500230020001E001B0019001600130010000D000A",
		INIT_79=>X"00200023002500270029002B002D002E002F002F0030003000300030002F002E",
		INIT_7A=>X"FFDFFFE4FFE8FFEDFFF1FFF6FFFAFFFF00030007000B000F00130017001A001D",
		INIT_7B=>X"FFAEFFAFFFB0FFB2FFB4FFB6FFB9FFBCFFBFFFC2FFC6FFCAFFCEFFD2FFD6FFDB",
		INIT_7C=>X"FFDDFFD7FFD1FFCBFFC6FFC2FFBDFFBAFFB7FFB4FFB2FFB0FFAFFFAEFFAEFFAE",
		INIT_7D=>X"0078006D00610056004B00400035002B00210017000E0005FFFCFFF4FFECFFE4",
		INIT_7E=>X"012A01200117010C010200F700ED00E100D600CB00BF00B300A7009C00900084",
		INIT_7F=>X"01780177017601750172016F016C01680163015E01580151014A0143013B0132",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_04,
		DOPADOP=>dopadop_04,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_05: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"0000000000FFFFFFFFFFFFFFFFFFFFFC0000000000000000000003FFFFFFFFFF",
		INITP_01=>X"FFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFF000000000000",
		INITP_02=>X"0000000FFFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFF",
		INITP_03=>X"FFFFFC0000000000000000000003FFFFFFFFFFFFFFFFFFFFFC00000000000000",
		INITP_04=>X"00003FFFFFFFFFFFFFFFFFFFFF0000000000000000000000FFFFFFFFFFFFFFFF",
		INITP_05=>X"FFF0000000000000000000000FFFFFFFFFFFFFFFFFFFFFC00000000000000000",
		INITP_06=>X"03FFFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFF",
		INITP_07=>X"0000000000000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000000000",
		INITP_08=>X"FFFFFFFFFFF000000000000000FFFFFFFFFFFFFFFC000000000000003FFFFFFF",
		INITP_09=>X"FFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFF0000000000000003FFFF",
		INITP_0A=>X"0FFFFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFF0000000000000003F",
		INITP_0B=>X"0000FFFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFF00000000000000",
		INITP_0C=>X"0000000FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFF00000000000",
		INITP_0D=>X"0000000000FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFC00000000",
		INITP_0E=>X"0000000000003FFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFFC00000",
		INITP_0F=>X"0000000000000003FFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFFC00",
		INIT_00=>X"FFFCFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_01=>X"00050004000400030003000200020001000100000000FFFFFFFEFFFEFFFDFFFD",
		INIT_02=>X"0007000700070007000800080007000700070007000700070006000600060005",
		INIT_03=>X"0000000100010002000300030004000400050005000500060006000600070007",
		INIT_04=>X"FFF8FFF9FFF9FFFAFFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFEFFFFFFFF0000",
		INIT_05=>X"FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF8",
		INIT_06=>X"0001000100000000FFFFFFFEFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFAFFF9",
		INIT_07=>X"0007000700070007000700060006000600050005000400040003000300020002",
		INIT_08=>X"0004000500050006000600060007000700070007000700080008000800080008",
		INIT_09=>X"FFFBFFFCFFFCFFFDFFFDFFFEFFFFFFFF00000000000100020002000300030004",
		INIT_0A=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFFAFFFAFFFB",
		INIT_0B=>X"FFFDFFFDFFFCFFFBFFFBFFFAFFFAFFFAFFF9FFF9FFF8FFF8FFF8FFF8FFF7FFF7",
		INIT_0C=>X"000600050005000500040004000300020002000100010000FFFFFFFFFFFEFFFE",
		INIT_0D=>X"0007000700080008000800080008000800080008000800070007000700070006",
		INIT_0E=>X"FFFF000000010001000200020003000300040004000500050006000600070007",
		INIT_0F=>X"FFF8FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFCFFFDFFFDFFFEFFFF",
		INIT_10=>X"FFF9FFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_11=>X"00020002000100010000FFFFFFFFFFFEFFFDFFFDFFFCFFFCFFFBFFFBFFFAFFFA",
		INIT_12=>X"0008000800080008000800080007000700070006000600050005000400040003",
		INIT_13=>X"0004000400050005000600060007000700070008000800080008000800080008",
		INIT_14=>X"FFFAFFFAFFFBFFFCFFFCFFFDFFFDFFFEFFFFFFFF000000010001000200030003",
		INIT_15=>X"FFF6FFF6FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9",
		INIT_16=>X"FFFEFFFDFFFDFFFCFFFBFFFBFFFAFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF7",
		INIT_17=>X"00080007000700060006000500040004000300030002000100010000FFFFFFFF",
		INIT_18=>X"0008000800080009000900090009000900090009000900090009000800080008",
		INIT_19=>X"FFFEFFFFFFFF0000000100020002000300040004000500050006000600070007",
		INIT_1A=>X"FFF6FFF6FFF6FFF7FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFD",
		INIT_1B=>X"FFF9FFF8FFF8FFF7FFF7FFF7FFF6FFF6FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF6",
		INIT_1C=>X"0004000400030002000100010000FFFFFFFEFFFEFFFDFFFCFFFBFFFBFFFAFFFA",
		INIT_1D=>X"000A000A000A000A000A000A0009000900090008000800070007000600060005",
		INIT_1E=>X"000300040005000600060007000700080008000900090009000A000A000A000A",
		INIT_1F=>X"FFF8FFF8FFF9FFF9FFFAFFFBFFFCFFFCFFFDFFFEFFFF00000000000100020003",
		INIT_20=>X"FFF5FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6FFF7",
		INIT_21=>X"FFFFFFFEFFFDFFFCFFFCFFFBFFFAFFF9FFF9FFF8FFF7FFF7FFF6FFF6FFF5FFF5",
		INIT_22=>X"000A000A00090009000800080007000600060005000400030002000100010000",
		INIT_23=>X"0009000A000A000B000B000B000C000C000C000C000C000C000C000B000B000B",
		INIT_24=>X"FFFCFFFDFFFEFFFF000000010002000200030004000500060007000700080009",
		INIT_25=>X"FFF2FFF2FFF3FFF3FFF3FFF4FFF4FFF5FFF6FFF6FFF7FFF8FFF9FFF9FFFAFFFB",
		INIT_26=>X"FFF8FFF7FFF6FFF6FFF5FFF5FFF4FFF4FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2",
		INIT_27=>X"000800070006000500040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9",
		INIT_28=>X"000E000E000E000E000E000E000E000D000D000D000C000B000B000A00090008",
		INIT_29=>X"0003000400050006000700080009000A000B000B000C000D000D000D000E000E",
		INIT_2A=>X"FFF3FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFBFFFDFFFEFFFF000000010002",
		INIT_2B=>X"FFF1FFF0FFF0FFEFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFF0FFF0FFF1FFF1FFF2",
		INIT_2C=>X"00010000FFFEFFFDFFFCFFFBFFF9FFF8FFF7FFF6FFF5FFF4FFF3FFF2FFF2FFF1",
		INIT_2D=>X"001100110010000F000E000E000D000C000B0009000800070006000500030002",
		INIT_2E=>X"000D000E000F0010001000110011001200120012001300130012001200120012",
		INIT_2F=>X"FFF7FFF9FFFAFFFCFFFDFFFF0000000200030005000600070009000A000B000C",
		INIT_30=>X"FFE9FFE9FFEAFFEAFFEBFFEBFFECFFEDFFEEFFEFFFF0FFF1FFF2FFF3FFF5FFF6",
		INIT_31=>X"FFF5FFF4FFF2FFF1FFF0FFEFFFEEFFEDFFECFFEBFFEBFFEAFFEAFFE9FFE9FFE9",
		INIT_32=>X"0010000F000D000B000A00080006000500030001FFFFFFFEFFFCFFFAFFF8FFF7",
		INIT_33=>X"001A001A001A001B001B001A001A001A00190018001700160015001400130012",
		INIT_34=>X"0003000500070009000B000D000F001000120013001500160017001800190019",
		INIT_35=>X"FFE3FFE5FFE6FFE8FFEAFFECFFEEFFF0FFF2FFF4FFF6FFF8FFFAFFFDFFFF0001",
		INIT_36=>X"FFE2FFE0FFDFFFDFFFDEFFDDFFDDFFDDFFDDFFDDFFDEFFDEFFDFFFE0FFE1FFE2",
		INIT_37=>X"000800050002FFFFFFFCFFF9FFF6FFF4FFF1FFEFFFECFFEAFFE8FFE6FFE5FFE3",
		INIT_38=>X"002D002C002A00290027002500230020001E001B0019001600130010000D000A",
		INIT_39=>X"00200023002500270029002B002D002E002F002F0030003000300030002F002E",
		INIT_3A=>X"FFDFFFE4FFE8FFEDFFF1FFF6FFFAFFFF00030007000B000F00130017001A001D",
		INIT_3B=>X"FFAEFFAFFFB0FFB2FFB4FFB6FFB9FFBCFFBFFFC2FFC6FFCAFFCEFFD2FFD6FFDB",
		INIT_3C=>X"FFDDFFD7FFD1FFCBFFC6FFC2FFBDFFBAFFB7FFB4FFB2FFB0FFAFFFAEFFAEFFAE",
		INIT_3D=>X"0078006D00610056004B00400035002B00210017000E0005FFFCFFF4FFECFFE4",
		INIT_3E=>X"012A01200117010C010200F700ED00E100D600CB00BF00B300A7009C00900084",
		INIT_3F=>X"01780177017601750172016F016C01680163015E01580151014A0143013B0132",
		INIT_40=>X"0000FFFFFFFEFFFEFFFDFFFCFFFBFFFBFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8",
		INIT_41=>X"0007000800070007000700070007000600060005000500040003000200020001",
		INIT_42=>X"FFFEFFFFFFFF0000000100020003000300040005000500060006000700070007",
		INIT_43=>X"FFF8FFF8FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFD",
		INIT_44=>X"0002000200010000FFFFFFFEFFFEFFFDFFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8",
		INIT_45=>X"0007000700070008000800080007000700070007000600060005000500040003",
		INIT_46=>X"FFFBFFFCFFFDFFFEFFFFFFFF0000000100020003000300040005000500060006",
		INIT_47=>X"FFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFB",
		INIT_48=>X"0005000400030002000200010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFFAFFF9",
		INIT_49=>X"0006000600070007000700080008000800080008000700070007000600060005",
		INIT_4A=>X"FFF9FFFAFFFBFFFCFFFCFFFDFFFEFFFF00000000000100020003000400040005",
		INIT_4B=>X"FFFAFFFAFFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9",
		INIT_4C=>X"0006000600050005000400030002000100010000FFFFFFFEFFFDFFFCFFFCFFFB",
		INIT_4D=>X"0004000500050006000600070007000800080008000800080008000800070007",
		INIT_4E=>X"FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFEFFFF00000001000100020003",
		INIT_4F=>X"FFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_50=>X"0008000700070007000600050005000400030002000100010000FFFFFFFEFFFD",
		INIT_51=>X"0002000300030004000500060006000700070008000800080008000800080008",
		INIT_52=>X"FFF7FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFEFFFF00000001",
		INIT_53=>X"FFFFFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_54=>X"0009000900080008000800070007000600060005000400030002000100000000",
		INIT_55=>X"FFFF000000010002000300040004000500060007000700080008000800090009",
		INIT_56=>X"FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFCFFFDFFFE",
		INIT_57=>X"00010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF6",
		INIT_58=>X"0009000900090009000900090009000800080007000700060005000400030002",
		INIT_59=>X"FFFCFFFDFFFEFFFF000000010002000300040005000600060007000800080009",
		INIT_5A=>X"FFF6FFF6FFF6FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF8FFF9FFF9FFFAFFFB",
		INIT_5B=>X"00040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF7FFF7",
		INIT_5C=>X"000800090009000A000A000A000A000A000A0009000900080008000700060005",
		INIT_5D=>X"FFF9FFFAFFFBFFFCFFFDFFFEFFFF000000010003000400050005000600070008",
		INIT_5E=>X"FFF7FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF7FFF7FFF8",
		INIT_5F=>X"00080007000600050004000300010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8",
		INIT_60=>X"0007000800090009000A000A000B000B000B000B000B000A000A000A00090008",
		INIT_61=>X"FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF000100020003000400050006",
		INIT_62=>X"FFF9FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF4FFF4FFF4FFF5FFF5",
		INIT_63=>X"000B000A000900080007000600050004000300010000FFFFFFFEFFFCFFFBFFFA",
		INIT_64=>X"00050006000700080009000A000B000B000C000C000C000C000C000C000C000B",
		INIT_65=>X"FFF3FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFCFFFDFFFE0000000100020004",
		INIT_66=>X"FFFCFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2",
		INIT_67=>X"000E000D000D000C000B000A00090008000700060004000300010000FFFFFFFD",
		INIT_68=>X"0001000300040006000700080009000A000B000C000D000D000E000E000E000E",
		INIT_69=>X"FFF0FFF0FFF1FFF1FFF2FFF3FFF3FFF5FFF6FFF7FFF8FFFAFFFBFFFDFFFE0000",
		INIT_6A=>X"0000FFFEFFFDFFFBFFF9FFF8FFF7FFF5FFF4FFF3FFF2FFF1FFF1FFF0FFF0FFF0",
		INIT_6B=>X"0010001000100010000F000F000E000D000C000B000900080006000500030002",
		INIT_6C=>X"FFFCFFFE000000020004000500070009000A000B000D000E000E000F00100010",
		INIT_6D=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEFFFF0FFF1FFF3FFF4FFF6FFF7FFF9FFFB",
		INIT_6E=>X"0006000400020000FFFEFFFCFFFAFFF8FFF6FFF5FFF3FFF2FFF0FFEFFFEFFFEE",
		INIT_6F=>X"00130013001400140014001400130013001200110010000E000D000B00090008",
		INIT_70=>X"FFF6FFF8FFFAFFFCFFFE00010003000500070009000B000D000E001000110012",
		INIT_71=>X"FFEBFFEAFFE9FFE9FFE8FFE8FFE8FFE9FFE9FFEAFFEBFFEDFFEEFFF0FFF2FFF3",
		INIT_72=>X"000E000C000A000700050002FFFFFFFDFFFAFFF8FFF6FFF4FFF1FFF0FFEEFFEC",
		INIT_73=>X"00150016001800190019001A001A001A001A0019001800170016001400120010",
		INIT_74=>X"FFEBFFEDFFF0FFF3FFF5FFF8FFFBFFFE000100040007000A000C000F00110013",
		INIT_75=>X"FFE9FFE7FFE5FFE4FFE2FFE1FFE0FFE0FFE0FFE0FFE1FFE2FFE3FFE5FFE7FFE9",
		INIT_76=>X"001C001A001700140010000D000A00060002FFFFFFFBFFF8FFF5FFF2FFEFFFEC",
		INIT_77=>X"00160019001C001F00210023002400250026002600260025002400220021001F",
		INIT_78=>X"FFD7FFDAFFDDFFE1FFE4FFE8FFEDFFF1FFF5FFFAFFFE00030007000B000F0013",
		INIT_79=>X"FFE8FFE4FFDFFFDBFFD8FFD5FFD3FFD1FFCFFFCFFFCEFFCFFFCFFFD0FFD2FFD4",
		INIT_7A=>X"003C003900350031002C00270021001B00160010000A0004FFFEFFF8FFF2FFED",
		INIT_7B=>X"0017001F0025002C00310036003A003E0041004300440044004400430042003F",
		INIT_7C=>X"FF95FF9AFFA0FFA7FFAEFFB6FFBFFFC8FFD1FFDAFFE3FFECFFF5FFFE0007000F",
		INIT_7D=>X"FFE8FFD8FFCAFFBEFFB3FFA9FFA1FF9AFF94FF90FF8DFF8BFF8BFF8CFF8EFF91",
		INIT_7E=>X"0145012E011600FE00E600CE00B6009F00870070005A00450030001C000AFFF8",
		INIT_7F=>X"021802170214020F0209020001F601EA01DD01CE01BE01AC019A01860171015B",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_05,
		DOPADOP=>dopadop_05,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_06: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFFFFFFFF000000000000000FFFFFFFFFFFFFFFC000000000000003FFFFFFF",
		INITP_01=>X"FFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFF0000000000000003FFFF",
		INITP_02=>X"0FFFFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFF0000000000000003F",
		INITP_03=>X"0000FFFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFF00000000000000",
		INITP_04=>X"0000000FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFF00000000000",
		INITP_05=>X"0000000000FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFC00000000",
		INITP_06=>X"0000000000003FFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFFC00000",
		INITP_07=>X"0000000000000003FFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFFC00",
		INITP_08=>X"FFFFF00000000003FFFFFFFFFFC00000000003FFFFFFFFFF00000000000FFFFF",
		INITP_09=>X"FFFFC0000000000FFFFFFFFFFF00000000003FFFFFFFFFFC0000000000FFFFFF",
		INITP_0A=>X"FFFC00000000003FFFFFFFFFF00000000000FFFFFFFFFFC00000000003FFFFFF",
		INITP_0B=>X"FFF00000000003FFFFFFFFFFC00000000003FFFFFFFFFF00000000000FFFFFFF",
		INITP_0C=>X"FFC0000000000FFFFFFFFFFF00000000003FFFFFFFFFFC0000000000FFFFFFFF",
		INITP_0D=>X"FC00000000003FFFFFFFFFF00000000000FFFFFFFFFFC00000000003FFFFFFFF",
		INITP_0E=>X"F00000000003FFFFFFFFFFC00000000003FFFFFFFFFF00000000000FFFFFFFFF",
		INITP_0F=>X"00000000000FFFFFFFFFFF00000000003FFFFFFFFFFC0000000000FFFFFFFFFF",
		INIT_00=>X"0000FFFFFFFEFFFEFFFDFFFCFFFBFFFBFFFAFFF9FFF9FFF9FFF8FFF8FFF8FFF8",
		INIT_01=>X"0007000800070007000700070007000600060005000500040003000200020001",
		INIT_02=>X"FFFEFFFFFFFF0000000100020003000300040005000500060006000700070007",
		INIT_03=>X"FFF8FFF8FFF7FFF7FFF8FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFBFFFBFFFCFFFD",
		INIT_04=>X"0002000200010000FFFFFFFEFFFEFFFDFFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8",
		INIT_05=>X"0007000700070008000800080007000700070007000600060005000500040003",
		INIT_06=>X"FFFBFFFCFFFDFFFEFFFFFFFF0000000100020003000300040005000500060006",
		INIT_07=>X"FFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9FFF9FFFAFFFAFFFB",
		INIT_08=>X"0005000400030002000200010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFFAFFF9",
		INIT_09=>X"0006000600070007000700080008000800080008000700070007000600060005",
		INIT_0A=>X"FFF9FFFAFFFBFFFCFFFCFFFDFFFEFFFF00000000000100020003000400040005",
		INIT_0B=>X"FFFAFFFAFFF9FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF8FFF8FFF9",
		INIT_0C=>X"0006000600050005000400030002000100010000FFFFFFFEFFFDFFFCFFFCFFFB",
		INIT_0D=>X"0004000500050006000600070007000800080008000800080008000800070007",
		INIT_0E=>X"FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFEFFFF00000001000100020003",
		INIT_0F=>X"FFFCFFFBFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_10=>X"0008000700070007000600050005000400030002000100010000FFFFFFFEFFFD",
		INIT_11=>X"0002000300030004000500060006000700070008000800080008000800080008",
		INIT_12=>X"FFF7FFF7FFF7FFF8FFF8FFF9FFF9FFFAFFFBFFFBFFFCFFFDFFFEFFFF00000001",
		INIT_13=>X"FFFFFFFEFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_14=>X"0009000900080008000800070007000600060005000400030002000100000000",
		INIT_15=>X"FFFF000000010002000300040004000500060007000700080008000800090009",
		INIT_16=>X"FFF6FFF6FFF6FFF6FFF6FFF7FFF7FFF8FFF8FFF9FFFAFFFAFFFBFFFCFFFDFFFE",
		INIT_17=>X"00010000FFFFFFFEFFFDFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF6",
		INIT_18=>X"0009000900090009000900090009000800080007000700060005000400030002",
		INIT_19=>X"FFFCFFFDFFFEFFFF000000010002000300040005000600060007000800080009",
		INIT_1A=>X"FFF6FFF6FFF6FFF5FFF5FFF5FFF6FFF6FFF6FFF7FFF7FFF8FFF9FFF9FFFAFFFB",
		INIT_1B=>X"00040003000200010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF7FFF7",
		INIT_1C=>X"000800090009000A000A000A000A000A000A0009000900080008000700060005",
		INIT_1D=>X"FFF9FFFAFFFBFFFCFFFDFFFEFFFF000000010003000400050005000600070008",
		INIT_1E=>X"FFF7FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF5FFF6FFF6FFF7FFF7FFF8",
		INIT_1F=>X"00080007000600050004000300010000FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8",
		INIT_20=>X"0007000800090009000A000A000B000B000B000B000B000A000A000A00090008",
		INIT_21=>X"FFF6FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF000100020003000400050006",
		INIT_22=>X"FFF9FFF8FFF7FFF6FFF5FFF5FFF4FFF4FFF4FFF3FFF3FFF4FFF4FFF4FFF5FFF5",
		INIT_23=>X"000B000A000900080007000600050004000300010000FFFFFFFEFFFCFFFBFFFA",
		INIT_24=>X"00050006000700080009000A000B000B000C000C000C000C000C000C000C000B",
		INIT_25=>X"FFF3FFF3FFF4FFF5FFF6FFF7FFF8FFF9FFFAFFFCFFFDFFFE0000000100020004",
		INIT_26=>X"FFFCFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF3FFF3FFF2FFF2FFF2FFF2FFF2FFF2",
		INIT_27=>X"000E000D000D000C000B000A00090008000700060004000300010000FFFFFFFD",
		INIT_28=>X"0001000300040006000700080009000A000B000C000D000D000E000E000E000E",
		INIT_29=>X"FFF0FFF0FFF1FFF1FFF2FFF3FFF3FFF5FFF6FFF7FFF8FFFAFFFBFFFDFFFE0000",
		INIT_2A=>X"0000FFFEFFFDFFFBFFF9FFF8FFF7FFF5FFF4FFF3FFF2FFF1FFF1FFF0FFF0FFF0",
		INIT_2B=>X"0010001000100010000F000F000E000D000C000B000900080006000500030002",
		INIT_2C=>X"FFFCFFFE000000020004000500070009000A000B000D000E000E000F00100010",
		INIT_2D=>X"FFEDFFEDFFEDFFEDFFEDFFEEFFEEFFEFFFF0FFF1FFF3FFF4FFF6FFF7FFF9FFFB",
		INIT_2E=>X"0006000400020000FFFEFFFCFFFAFFF8FFF6FFF5FFF3FFF2FFF0FFEFFFEFFFEE",
		INIT_2F=>X"00130013001400140014001400130013001200110010000E000D000B00090008",
		INIT_30=>X"FFF6FFF8FFFAFFFCFFFE00010003000500070009000B000D000E001000110012",
		INIT_31=>X"FFEBFFEAFFE9FFE9FFE8FFE8FFE8FFE9FFE9FFEAFFEBFFEDFFEEFFF0FFF2FFF3",
		INIT_32=>X"000E000C000A000700050002FFFFFFFDFFFAFFF8FFF6FFF4FFF1FFF0FFEEFFEC",
		INIT_33=>X"00150016001800190019001A001A001A001A0019001800170016001400120010",
		INIT_34=>X"FFEBFFEDFFF0FFF3FFF5FFF8FFFBFFFE000100040007000A000C000F00110013",
		INIT_35=>X"FFE9FFE7FFE5FFE4FFE2FFE1FFE0FFE0FFE0FFE0FFE1FFE2FFE3FFE5FFE7FFE9",
		INIT_36=>X"001C001A001700140010000D000A00060002FFFFFFFBFFF8FFF5FFF2FFEFFFEC",
		INIT_37=>X"00160019001C001F00210023002400250026002600260025002400220021001F",
		INIT_38=>X"FFD7FFDAFFDDFFE1FFE4FFE8FFEDFFF1FFF5FFFAFFFE00030007000B000F0013",
		INIT_39=>X"FFE8FFE4FFDFFFDBFFD8FFD5FFD3FFD1FFCFFFCFFFCEFFCFFFCFFFD0FFD2FFD4",
		INIT_3A=>X"003C003900350031002C00270021001B00160010000A0004FFFEFFF8FFF2FFED",
		INIT_3B=>X"0017001F0025002C00310036003A003E0041004300440044004400430042003F",
		INIT_3C=>X"FF95FF9AFFA0FFA7FFAEFFB6FFBFFFC8FFD1FFDAFFE3FFECFFF5FFFE0007000F",
		INIT_3D=>X"FFE8FFD8FFCAFFBEFFB3FFA9FFA1FF9AFF94FF90FF8DFF8BFF8BFF8CFF8EFF91",
		INIT_3E=>X"0145012E011600FE00E600CE00B6009F00870070005A00450030001C000AFFF8",
		INIT_3F=>X"021802170214020F0209020001F601EA01DD01CE01BE01AC019A01860171015B",
		INIT_40=>X"000500040003000200010000FFFFFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8FFF8",
		INIT_41=>X"0000000100020003000400050006000700070007000700070007000700060006",
		INIT_42=>X"FFF9FFF9FFF8FFF8FFF8FFF7FFF8FFF8FFF8FFF9FFFAFFFAFFFBFFFCFFFEFFFF",
		INIT_43=>X"00070007000700060006000500040003000200010000FFFEFFFDFFFCFFFBFFFA",
		INIT_44=>X"FFFBFFFCFFFDFFFEFFFF00000001000200030004000500060007000700070008",
		INIT_45=>X"FFFEFFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF8FFF8FFF8FFF9FFFA",
		INIT_46=>X"000600070007000700080008000700070006000600050004000300020001FFFF",
		INIT_47=>X"FFF8FFF8FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF000000010002000400050005",
		INIT_48=>X"0004000300020001FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF8FFF7FFF7",
		INIT_49=>X"0002000300040005000600060007000700080008000800070007000600060005",
		INIT_4A=>X"FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF0000",
		INIT_4B=>X"000800070006000600050004000300020000FFFFFFFEFFFDFFFCFFFBFFFAFFF9",
		INIT_4C=>X"FFFCFFFDFFFEFFFF000000020003000400050006000700070008000800080008",
		INIT_4D=>X"FFFDFFFCFFFAFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFB",
		INIT_4E=>X"00070008000800080008000800070007000600050004000300020000FFFFFFFE",
		INIT_4F=>X"FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF0001000200030004000500060007",
		INIT_50=>X"000300010000FFFFFFFEFFFCFFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7",
		INIT_51=>X"0003000400050006000700080008000800080008000800070007000600050004",
		INIT_52=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFE000000010002",
		INIT_53=>X"00070007000600050004000300010000FFFFFFFDFFFCFFFBFFFAFFF9FFF8FFF7",
		INIT_54=>X"FFFDFFFE00000001000200040005000600070007000800080009000900080008",
		INIT_55=>X"FFFBFFFAFFF9FFF8FFF7FFF7FFF6FFF6FFF6FFF7FFF7FFF8FFF9FFFAFFFBFFFC",
		INIT_56=>X"0009000900090009000800080007000600050004000300010000FFFFFFFDFFFC",
		INIT_57=>X"FFF7FFF8FFF9FFFBFFFCFFFDFFFE000000010003000400050006000700080008",
		INIT_58=>X"00010000FFFEFFFDFFFCFFFAFFF9FFF8FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF7",
		INIT_59=>X"0005000700070008000900090009000900090009000800070006000500040003",
		INIT_5A=>X"FFF5FFF5FFF6FFF6FFF6FFF7FFF8FFF9FFFAFFFCFFFDFFFF0000000100030004",
		INIT_5B=>X"0008000600050004000300010000FFFEFFFDFFFBFFFAFFF9FFF8FFF7FFF6FFF6",
		INIT_5C=>X"FFFF000000020003000500060007000800090009000A000A000A000A00090008",
		INIT_5D=>X"FFF8FFF7FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF6FFF7FFF8FFF9FFFAFFFCFFFD",
		INIT_5E=>X"000B000A000A000A0009000800070005000400030001FFFFFFFEFFFCFFFBFFF9",
		INIT_5F=>X"FFF8FFF9FFFAFFFCFFFDFFFF00000002000400050006000800090009000A000A",
		INIT_60=>X"FFFFFFFEFFFCFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF4FFF4FFF4FFF5FFF6FFF6",
		INIT_61=>X"00080009000A000B000B000B000B000B000A0009000800070006000400030001",
		INIT_62=>X"FFF3FFF4FFF4FFF5FFF6FFF7FFF8FFFAFFFCFFFDFFFF00010002000400060007",
		INIT_63=>X"00070006000400030001FFFFFFFDFFFBFFFAFFF8FFF7FFF6FFF5FFF4FFF3FFF3",
		INIT_64=>X"000100030005000600080009000A000B000C000C000C000C000C000B000A0009",
		INIT_65=>X"FFF5FFF4FFF3FFF2FFF2FFF2FFF3FFF3FFF4FFF5FFF7FFF8FFFAFFFBFFFDFFFF",
		INIT_66=>X"000D000D000C000B000A00080006000500030001FFFFFFFDFFFBFFF9FFF7FFF6",
		INIT_67=>X"FFF8FFF9FFFBFFFDFFFF00010003000500070009000A000B000C000D000D000D",
		INIT_68=>X"FFFCFFFAFFF8FFF6FFF5FFF3FFF2FFF2FFF1FFF1FFF1FFF1FFF2FFF3FFF4FFF6",
		INIT_69=>X"000D000E000F000F000F000F000E000D000C000A00090007000500030001FFFE",
		INIT_6A=>X"FFF0FFF1FFF2FFF3FFF5FFF7FFF9FFFBFFFD00000002000400060008000A000C",
		INIT_6B=>X"0008000500030000FFFEFFFCFFF9FFF7FFF5FFF3FFF2FFF1FFF0FFEFFFEFFFEF",
		INIT_6C=>X"00050007000A000C000D000F001000100011001100100010000F000D000C000A",
		INIT_6D=>X"FFEFFFEEFFEDFFEDFFEDFFEEFFEFFFF0FFF2FFF4FFF6FFF8FFFBFFFD00000003",
		INIT_6E=>X"00120011000F000D000B0008000600030000FFFDFFFBFFF8FFF6FFF3FFF2FFF0",
		INIT_6F=>X"FFF8FFFAFFFD0000000300060009000B000E0010001100120013001300130013",
		INIT_70=>X"FFF6FFF4FFF1FFEFFFEDFFECFFEBFFEAFFEAFFEAFFEBFFECFFEEFFF0FFF2FFF5",
		INIT_71=>X"00160017001700170016001500130011000F000C000A000600030000FFFDFFFA",
		INIT_72=>X"FFE9FFEBFFEDFFF0FFF3FFF6FFFAFFFD000100050008000B000E001100130015",
		INIT_73=>X"000700040000FFFCFFF8FFF4FFF1FFEEFFEBFFE9FFE7FFE6FFE6FFE6FFE6FFE7",
		INIT_74=>X"000E001200150018001A001B001C001C001C001B001A001800150012000F000B",
		INIT_75=>X"FFE0FFDFFFDFFFE0FFE1FFE3FFE6FFE9FFECFFF0FFF5FFF9FFFD00020006000A",
		INIT_76=>X"001E001B00170013000E00090004FFFFFFFAFFF5FFF1FFECFFE9FFE5FFE3FFE1",
		INIT_77=>X"FFF7FFFD00030009000E00140018001C001F0022002400250025002400230021",
		INIT_78=>X"FFE5FFE0FFDBFFD8FFD5FFD4FFD3FFD4FFD5FFD7FFDAFFDDFFE2FFE7FFECFFF2",
		INIT_79=>X"0035003500340032002F002B00260020001A0013000C0005FFFEFFF7FFF0FFEA",
		INIT_7A=>X"FFCCFFD3FFDBFFE3FFECFFF5FFFD0006000F0017001E0024002A002E00320034",
		INIT_7B=>X"0008FFFCFFF0FFE6FFDCFFD3FFCBFFC5FFC0FFBCFFBAFFBAFFBBFFBDFFC1FFC6",
		INIT_7C=>X"004700500058005D006000610060005D00580052004A00410036002B001F0014",
		INIT_7D=>X"FF5DFF62FF6BFF76FF83FF92FFA2FFB4FFC6FFD9FFEBFFFD000F001F002E003B",
		INIT_7E=>X"00EC00BD008F0063003A0014FFF0FFD0FFB4FF9BFF87FF76FF69FF60FF5CFF5A",
		INIT_7F=>X"02F802F502ED02E002CD02B6029A027A02570230020601D901AB017C014C011B",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_06,
		DOPADOP=>dopadop_06,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_07: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFF00000000003FFFFFFFFFFC00000000003FFFFFFFFFF00000000000FFFFF",
		INITP_01=>X"FFFFC0000000000FFFFFFFFFFF00000000003FFFFFFFFFFC0000000000FFFFFF",
		INITP_02=>X"FFFC00000000003FFFFFFFFFF00000000000FFFFFFFFFFC00000000003FFFFFF",
		INITP_03=>X"FFF00000000003FFFFFFFFFFC00000000003FFFFFFFFFF00000000000FFFFFFF",
		INITP_04=>X"FFC0000000000FFFFFFFFFFF00000000003FFFFFFFFFFC0000000000FFFFFFFF",
		INITP_05=>X"FC00000000003FFFFFFFFFF00000000000FFFFFFFFFFC00000000003FFFFFFFF",
		INITP_06=>X"F00000000003FFFFFFFFFFC00000000003FFFFFFFFFF00000000000FFFFFFFFF",
		INITP_07=>X"00000000000FFFFFFFFFFF00000000003FFFFFFFFFFC0000000000FFFFFFFFFF",
		INITP_08=>X"FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC00000003FFFFFFF00000003FFF",
		INITP_09=>X"000FFFFFFFC00000003FFFFFFF00000003FFFFFFF00000003FFFFFFF00000000",
		INITP_0A=>X"0000003FFFFFFF00000003FFFFFFF00000000FFFFFFFC0000000FFFFFFFC0000",
		INITP_0B=>X"FF00000003FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFF0",
		INITP_0C=>X"FFFFFC0000000FFFFFFFC0000000FFFFFFFF00000003FFFFFFF00000003FFFFF",
		INITP_0D=>X"0FFFFFFFF00000003FFFFFFF00000003FFFFFFF00000003FFFFFFFC0000000FF",
		INITP_0E=>X"00003FFFFFFF00000003FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC000000",
		INITP_0F=>X"00000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFF00000003FFFFFFF000",
		INIT_00=>X"000500040003000200010000FFFFFFFDFFFCFFFBFFFAFFFAFFF9FFF8FFF8FFF8",
		INIT_01=>X"0000000100020003000400050006000700070007000700070007000700060006",
		INIT_02=>X"FFF9FFF9FFF8FFF8FFF8FFF7FFF8FFF8FFF8FFF9FFFAFFFAFFFBFFFCFFFEFFFF",
		INIT_03=>X"00070007000700060006000500040003000200010000FFFEFFFDFFFCFFFBFFFA",
		INIT_04=>X"FFFBFFFCFFFDFFFEFFFF00000001000200030004000500060007000700070008",
		INIT_05=>X"FFFEFFFDFFFCFFFBFFFAFFF9FFF9FFF8FFF8FFF7FFF7FFF8FFF8FFF8FFF9FFFA",
		INIT_06=>X"000600070007000700080008000700070006000600050004000300020001FFFF",
		INIT_07=>X"FFF8FFF8FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF000000010002000400050005",
		INIT_08=>X"0004000300020001FFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF8FFF8FFF7FFF7",
		INIT_09=>X"0002000300040005000600060007000700080008000800070007000600060005",
		INIT_0A=>X"FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF0000",
		INIT_0B=>X"000800070006000600050004000300020000FFFFFFFEFFFDFFFCFFFBFFFAFFF9",
		INIT_0C=>X"FFFCFFFDFFFEFFFF000000020003000400050006000700070008000800080008",
		INIT_0D=>X"FFFDFFFCFFFAFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF8FFF8FFF9FFFAFFFB",
		INIT_0E=>X"00070008000800080008000800070007000600050004000300020000FFFFFFFE",
		INIT_0F=>X"FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFEFFFF0001000200030004000500060007",
		INIT_10=>X"000300010000FFFFFFFEFFFCFFFBFFFAFFF9FFF8FFF8FFF7FFF7FFF7FFF7FFF7",
		INIT_11=>X"0003000400050006000700080008000800080008000800070007000600050004",
		INIT_12=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF8FFF9FFFAFFFBFFFCFFFDFFFE000000010002",
		INIT_13=>X"00070007000600050004000300010000FFFFFFFDFFFCFFFBFFFAFFF9FFF8FFF7",
		INIT_14=>X"FFFDFFFE00000001000200040005000600070007000800080009000900080008",
		INIT_15=>X"FFFBFFFAFFF9FFF8FFF7FFF7FFF6FFF6FFF6FFF7FFF7FFF8FFF9FFFAFFFBFFFC",
		INIT_16=>X"0009000900090009000800080007000600050004000300010000FFFFFFFDFFFC",
		INIT_17=>X"FFF7FFF8FFF9FFFBFFFCFFFDFFFE000000010003000400050006000700080008",
		INIT_18=>X"00010000FFFEFFFDFFFCFFFAFFF9FFF8FFF7FFF7FFF6FFF6FFF6FFF6FFF6FFF7",
		INIT_19=>X"0005000700070008000900090009000900090009000800070006000500040003",
		INIT_1A=>X"FFF5FFF5FFF6FFF6FFF6FFF7FFF8FFF9FFFAFFFCFFFDFFFF0000000100030004",
		INIT_1B=>X"0008000600050004000300010000FFFEFFFDFFFBFFFAFFF9FFF8FFF7FFF6FFF6",
		INIT_1C=>X"FFFF000000020003000500060007000800090009000A000A000A000A00090008",
		INIT_1D=>X"FFF8FFF7FFF6FFF6FFF5FFF5FFF5FFF5FFF5FFF6FFF7FFF8FFF9FFFAFFFCFFFD",
		INIT_1E=>X"000B000A000A000A0009000800070005000400030001FFFFFFFEFFFCFFFBFFF9",
		INIT_1F=>X"FFF8FFF9FFFAFFFCFFFDFFFF00000002000400050006000800090009000A000A",
		INIT_20=>X"FFFFFFFEFFFCFFFAFFF9FFF8FFF7FFF6FFF5FFF4FFF4FFF4FFF4FFF5FFF6FFF6",
		INIT_21=>X"00080009000A000B000B000B000B000B000A0009000800070006000400030001",
		INIT_22=>X"FFF3FFF4FFF4FFF5FFF6FFF7FFF8FFFAFFFCFFFDFFFF00010002000400060007",
		INIT_23=>X"00070006000400030001FFFFFFFDFFFBFFFAFFF8FFF7FFF6FFF5FFF4FFF3FFF3",
		INIT_24=>X"000100030005000600080009000A000B000C000C000C000C000C000B000A0009",
		INIT_25=>X"FFF5FFF4FFF3FFF2FFF2FFF2FFF3FFF3FFF4FFF5FFF7FFF8FFFAFFFBFFFDFFFF",
		INIT_26=>X"000D000D000C000B000A00080006000500030001FFFFFFFDFFFBFFF9FFF7FFF6",
		INIT_27=>X"FFF8FFF9FFFBFFFDFFFF00010003000500070009000A000B000C000D000D000D",
		INIT_28=>X"FFFCFFFAFFF8FFF6FFF5FFF3FFF2FFF2FFF1FFF1FFF1FFF1FFF2FFF3FFF4FFF6",
		INIT_29=>X"000D000E000F000F000F000F000E000D000C000A00090007000500030001FFFE",
		INIT_2A=>X"FFF0FFF1FFF2FFF3FFF5FFF7FFF9FFFBFFFD00000002000400060008000A000C",
		INIT_2B=>X"0008000500030000FFFEFFFCFFF9FFF7FFF5FFF3FFF2FFF1FFF0FFEFFFEFFFEF",
		INIT_2C=>X"00050007000A000C000D000F001000100011001100100010000F000D000C000A",
		INIT_2D=>X"FFEFFFEEFFEDFFEDFFEDFFEEFFEFFFF0FFF2FFF4FFF6FFF8FFFBFFFD00000003",
		INIT_2E=>X"00120011000F000D000B0008000600030000FFFDFFFBFFF8FFF6FFF3FFF2FFF0",
		INIT_2F=>X"FFF8FFFAFFFD0000000300060009000B000E0010001100120013001300130013",
		INIT_30=>X"FFF6FFF4FFF1FFEFFFEDFFECFFEBFFEAFFEAFFEAFFEBFFECFFEEFFF0FFF2FFF5",
		INIT_31=>X"00160017001700170016001500130011000F000C000A000600030000FFFDFFFA",
		INIT_32=>X"FFE9FFEBFFEDFFF0FFF3FFF6FFFAFFFD000100050008000B000E001100130015",
		INIT_33=>X"000700040000FFFCFFF8FFF4FFF1FFEEFFEBFFE9FFE7FFE6FFE6FFE6FFE6FFE7",
		INIT_34=>X"000E001200150018001A001B001C001C001C001B001A001800150012000F000B",
		INIT_35=>X"FFE0FFDFFFDFFFE0FFE1FFE3FFE6FFE9FFECFFF0FFF5FFF9FFFD00020006000A",
		INIT_36=>X"001E001B00170013000E00090004FFFFFFFAFFF5FFF1FFECFFE9FFE5FFE3FFE1",
		INIT_37=>X"FFF7FFFD00030009000E00140018001C001F0022002400250025002400230021",
		INIT_38=>X"FFE5FFE0FFDBFFD8FFD5FFD4FFD3FFD4FFD5FFD7FFDAFFDDFFE2FFE7FFECFFF2",
		INIT_39=>X"0035003500340032002F002B00260020001A0013000C0005FFFEFFF7FFF0FFEA",
		INIT_3A=>X"FFCCFFD3FFDBFFE3FFECFFF5FFFD0006000F0017001E0024002A002E00320034",
		INIT_3B=>X"0008FFFCFFF0FFE6FFDCFFD3FFCBFFC5FFC0FFBCFFBAFFBAFFBBFFBDFFC1FFC6",
		INIT_3C=>X"004700500058005D006000610060005D00580052004A00410036002B001F0014",
		INIT_3D=>X"FF5DFF62FF6BFF76FF83FF92FFA2FFB4FFC6FFD9FFEBFFFD000F001F002E003B",
		INIT_3E=>X"00EC00BD008F0063003A0014FFF0FFD0FFB4FF9BFF87FF76FF69FF60FF5CFF5A",
		INIT_3F=>X"02F802F502ED02E002CD02B6029A027A02570230020601D901AB017C014C011B",
		INIT_40=>X"000700070007000700060005000300020000FFFFFFFDFFFBFFFAFFF9FFF8FFF8",
		INIT_41=>X"FFF8FFF8FFF8FFF8FFF8FFF9FFFBFFFCFFFDFFFF000100020004000500060007",
		INIT_42=>X"00060007000700070007000600050004000300010000FFFEFFFCFFFBFFFAFFF9",
		INIT_43=>X"FFF9FFF8FFF8FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFE00000001000300040006",
		INIT_44=>X"000500060007000700080007000700060005000400020001FFFFFFFDFFFCFFFA",
		INIT_45=>X"FFFBFFFAFFF9FFF8FFF8FFF7FFF8FFF8FFF9FFFAFFFBFFFDFFFF000000020003",
		INIT_46=>X"00020004000500060007000700080007000700060005000300020000FFFEFFFD",
		INIT_47=>X"FFFEFFFCFFFBFFFAFFF9FFF8FFF7FFF7FFF8FFF8FFF9FFFAFFFCFFFDFFFF0001",
		INIT_48=>X"0000000100030004000600070007000800080007000700060004000300010000",
		INIT_49=>X"0001FFFFFFFDFFFCFFFAFFF9FFF8FFF8FFF7FFF7FFF8FFF9FFFAFFFBFFFCFFFE",
		INIT_4A=>X"FFFDFFFF00000002000400050006000700080008000800070006000500040002",
		INIT_4B=>X"000300020000FFFEFFFDFFFBFFFAFFF9FFF8FFF7FFF7FFF7FFF8FFF9FFFAFFFB",
		INIT_4C=>X"FFFAFFFCFFFDFFFF000100030004000500070007000800080008000700060005",
		INIT_4D=>X"00060004000300010000FFFEFFFCFFFBFFF9FFF8FFF8FFF7FFF7FFF7FFF8FFF9",
		INIT_4E=>X"FFF8FFF9FFFBFFFCFFFE00000001000300050006000700080008000800080007",
		INIT_4F=>X"000800070005000400020001FFFFFFFDFFFCFFFAFFF9FFF8FFF7FFF7FFF7FFF7",
		INIT_50=>X"FFF7FFF8FFF8FFFAFFFBFFFDFFFF000000020004000500060007000800080008",
		INIT_51=>X"00080008000700060005000400020000FFFEFFFDFFFBFFF9FFF8FFF7FFF7FFF7",
		INIT_52=>X"FFF7FFF7FFF7FFF8FFF9FFFAFFFCFFFDFFFF0001000300040006000700080008",
		INIT_53=>X"0008000900080008000700060005000300010000FFFEFFFCFFFAFFF9FFF8FFF7",
		INIT_54=>X"FFF7FFF7FFF6FFF6FFF7FFF8FFF9FFFAFFFCFFFE000000020003000500060007",
		INIT_55=>X"00070008000900090009000800070006000400030001FFFFFFFDFFFBFFFAFFF8",
		INIT_56=>X"FFF9FFF8FFF7FFF6FFF6FFF6FFF7FFF8FFF9FFFBFFFDFFFF0000000200040006",
		INIT_57=>X"0005000600080008000900090009000800070006000400020000FFFEFFFCFFFB",
		INIT_58=>X"FFFCFFFAFFF8FFF7FFF6FFF6FFF6FFF6FFF7FFF8FFFAFFFBFFFDFFFF00010003",
		INIT_59=>X"00020004000600070008000900090009000900080007000500030001FFFFFFFD",
		INIT_5A=>X"FFFFFFFDFFFBFFF9FFF8FFF6FFF6FFF5FFF6FFF6FFF7FFF8FFFAFFFCFFFE0000",
		INIT_5B=>X"FFFE000100030005000600080009000A000A000A000900080006000500030001",
		INIT_5C=>X"00020000FFFEFFFCFFFAFFF8FFF7FFF6FFF5FFF5FFF5FFF6FFF7FFF9FFFAFFFC",
		INIT_5D=>X"FFFBFFFDFFFF00010004000500070009000A000A000A000A0009000800060004",
		INIT_5E=>X"000600040002FFFFFFFDFFFBFFF9FFF7FFF6FFF5FFF5FFF5FFF5FFF6FFF7FFF9",
		INIT_5F=>X"FFF8FFF9FFFBFFFE000000020004000600080009000A000B000B000A00090008",
		INIT_60=>X"00090007000500030001FFFFFFFCFFFAFFF8FFF6FFF5FFF4FFF4FFF4FFF5FFF6",
		INIT_61=>X"FFF5FFF6FFF8FFFAFFFCFFFE00010003000500070009000A000B000B000B000A",
		INIT_62=>X"000B000A00090007000500030000FFFEFFFBFFF9FFF7FFF6FFF4FFF4FFF4FFF4",
		INIT_63=>X"FFF3FFF3FFF5FFF6FFF8FFFAFFFDFFFF0002000400060008000A000B000C000C",
		INIT_64=>X"000C000C000C000B0009000700050002FFFFFFFDFFFAFFF8FFF6FFF5FFF3FFF3",
		INIT_65=>X"FFF2FFF2FFF2FFF3FFF4FFF6FFF8FFFBFFFD0000000300050008000A000B000C",
		INIT_66=>X"000C000D000D000D000C000B0009000700040001FFFEFFFCFFF9FFF7FFF5FFF3",
		INIT_67=>X"FFF4FFF2FFF1FFF1FFF2FFF3FFF4FFF6FFF9FFFBFFFE0001000400070009000B",
		INIT_68=>X"000A000C000D000E000E000E000D000B0009000600030000FFFDFFFAFFF8FFF5",
		INIT_69=>X"FFF6FFF4FFF2FFF1FFF0FFF0FFF1FFF2FFF4FFF6FFF9FFFCFFFF000200050008",
		INIT_6A=>X"0007000A000C000E000F000F000F000E000D000B000800060002FFFFFFFCFFF9",
		INIT_6B=>X"FFFBFFF7FFF5FFF2FFF0FFEFFFEFFFEFFFF0FFF2FFF4FFF7FFFAFFFD00000004",
		INIT_6C=>X"000200050009000B000E0010001100110010000F000E000B000800050002FFFE",
		INIT_6D=>X"0000FFFDFFF9FFF5FFF3FFF0FFEEFFEDFFEDFFEEFFEFFFF1FFF4FFF7FFFAFFFE",
		INIT_6E=>X"FFFBFFFF00030007000B000E001000120013001300120010000E000B00080004",
		INIT_6F=>X"00080003FFFFFFFBFFF7FFF3FFF0FFEEFFECFFEBFFEBFFECFFEEFFF1FFF4FFF7",
		INIT_70=>X"FFF4FFF8FFFC000100050009000D0010001300140015001500130011000F000B",
		INIT_71=>X"000F000B00070002FFFDFFF9FFF4FFF0FFEDFFEBFFE9FFE9FFE9FFEBFFEDFFF0",
		INIT_72=>X"FFEBFFEFFFF4FFF8FFFE00030008000C00100013001600170018001700150013",
		INIT_73=>X"001800150010000C00060001FFFBFFF6FFF1FFEDFFEAFFE7FFE6FFE6FFE7FFE8",
		INIT_74=>X"FFE3FFE6FFE9FFEEFFF3FFF9FFFF0005000B001000140018001A001B001B001A",
		INIT_75=>X"0020001E001B00170012000C0005FFFFFFF8FFF2FFEDFFE8FFE5FFE2FFE1FFE2",
		INIT_76=>X"FFDBFFDCFFDEFFE2FFE7FFEDFFF3FFFA00020009000F0015001A001D00200021",
		INIT_77=>X"00280028002700240020001A0013000C0004FFFCFFF4FFEDFFE7FFE2FFDEFFDC",
		INIT_78=>X"FFD4FFD2FFD2FFD3FFD7FFDCFFE3FFEBFFF3FFFC0005000E0015001C00220026",
		INIT_79=>X"002E0033003400340032002D0027001F0016000C0001FFF7FFEEFFE5FFDEFFD8",
		INIT_7A=>X"FFCEFFC7FFC3FFC1FFC2FFC5FFCBFFD3FFDDFFE8FFF3FFFF000B001600200028",
		INIT_7B=>X"0033003E0046004B004C004A0045003E00330027001A000CFFFDFFF0FFE3FFD7",
		INIT_7C=>X"FFCAFFB9FFACFFA3FF9EFF9DFFA1FFA8FFB3FFC0FFD0FFE1FFF3000500160026",
		INIT_7D=>X"003600520069007A0085008A00890082007600660052003C0024000CFFF4FFDE",
		INIT_7E=>X"FFC8FF8EFF5FFF3CFF24FF17FF15FF1DFF2DFF45FF62FF84FFA9FFCEFFF30016",
		INIT_7F=>X"04380430041903F303C00381033602E30289022A01C90168010900AE0059000C",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_07,
		DOPADOP=>dopadop_07,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_08: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC00000003FFFFFFF00000003FFF",
		INITP_01=>X"000FFFFFFFC00000003FFFFFFF00000003FFFFFFF00000003FFFFFFF00000000",
		INITP_02=>X"0000003FFFFFFF00000003FFFFFFF00000000FFFFFFFC0000000FFFFFFFC0000",
		INITP_03=>X"FF00000003FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFF0",
		INITP_04=>X"FFFFFC0000000FFFFFFFC0000000FFFFFFFF00000003FFFFFFF00000003FFFFF",
		INITP_05=>X"0FFFFFFFF00000003FFFFFFF00000003FFFFFFF00000003FFFFFFFC0000000FF",
		INITP_06=>X"00003FFFFFFF00000003FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC000000",
		INITP_07=>X"00000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFF00000003FFFFFFF000",
		INITP_08=>X"00FFFFFC00000FFFFF000003FFFFF000003FFFFF000003FFFFC00000FFFFFC00",
		INITP_09=>X"0FFFFFC00000FFFFF000003FFFFF000003FFFFF000003FFFFC00000FFFFFC000",
		INITP_0A=>X"FFFFFC00003FFFFF000003FFFFF000003FFFFF000003FFFFC00000FFFFFC0000",
		INITP_0B=>X"FFFFC00003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000",
		INITP_0C=>X"FFFC00003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000F",
		INITP_0D=>X"FFC00003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000FF",
		INITP_0E=>X"FC00003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000FFF",
		INITP_0F=>X"000003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000FFFF",
		INIT_00=>X"000700070007000700060005000300020000FFFFFFFDFFFBFFFAFFF9FFF8FFF8",
		INIT_01=>X"FFF8FFF8FFF8FFF8FFF8FFF9FFFBFFFCFFFDFFFF000100020004000500060007",
		INIT_02=>X"00060007000700070007000600050004000300010000FFFEFFFCFFFBFFFAFFF9",
		INIT_03=>X"FFF9FFF8FFF8FFF7FFF8FFF8FFF9FFFAFFFBFFFCFFFE00000001000300040006",
		INIT_04=>X"000500060007000700080007000700060005000400020001FFFFFFFDFFFCFFFA",
		INIT_05=>X"FFFBFFFAFFF9FFF8FFF8FFF7FFF8FFF8FFF9FFFAFFFBFFFDFFFF000000020003",
		INIT_06=>X"00020004000500060007000700080007000700060005000300020000FFFEFFFD",
		INIT_07=>X"FFFEFFFCFFFBFFFAFFF9FFF8FFF7FFF7FFF8FFF8FFF9FFFAFFFCFFFDFFFF0001",
		INIT_08=>X"0000000100030004000600070007000800080007000700060004000300010000",
		INIT_09=>X"0001FFFFFFFDFFFCFFFAFFF9FFF8FFF8FFF7FFF7FFF8FFF9FFFAFFFBFFFCFFFE",
		INIT_0A=>X"FFFDFFFF00000002000400050006000700080008000800070006000500040002",
		INIT_0B=>X"000300020000FFFEFFFDFFFBFFFAFFF9FFF8FFF7FFF7FFF7FFF8FFF9FFFAFFFB",
		INIT_0C=>X"FFFAFFFCFFFDFFFF000100030004000500070007000800080008000700060005",
		INIT_0D=>X"00060004000300010000FFFEFFFCFFFBFFF9FFF8FFF8FFF7FFF7FFF7FFF8FFF9",
		INIT_0E=>X"FFF8FFF9FFFBFFFCFFFE00000001000300050006000700080008000800080007",
		INIT_0F=>X"000800070005000400020001FFFFFFFDFFFCFFFAFFF9FFF8FFF7FFF7FFF7FFF7",
		INIT_10=>X"FFF7FFF8FFF8FFFAFFFBFFFDFFFF000000020004000500060007000800080008",
		INIT_11=>X"00080008000700060005000400020000FFFEFFFDFFFBFFF9FFF8FFF7FFF7FFF7",
		INIT_12=>X"FFF7FFF7FFF7FFF8FFF9FFFAFFFCFFFDFFFF0001000300040006000700080008",
		INIT_13=>X"0008000900080008000700060005000300010000FFFEFFFCFFFAFFF9FFF8FFF7",
		INIT_14=>X"FFF7FFF7FFF6FFF6FFF7FFF8FFF9FFFAFFFCFFFE000000020003000500060007",
		INIT_15=>X"00070008000900090009000800070006000400030001FFFFFFFDFFFBFFFAFFF8",
		INIT_16=>X"FFF9FFF8FFF7FFF6FFF6FFF6FFF7FFF8FFF9FFFBFFFDFFFF0000000200040006",
		INIT_17=>X"0005000600080008000900090009000800070006000400020000FFFEFFFCFFFB",
		INIT_18=>X"FFFCFFFAFFF8FFF7FFF6FFF6FFF6FFF6FFF7FFF8FFFAFFFBFFFDFFFF00010003",
		INIT_19=>X"00020004000600070008000900090009000900080007000500030001FFFFFFFD",
		INIT_1A=>X"FFFFFFFDFFFBFFF9FFF8FFF6FFF6FFF5FFF6FFF6FFF7FFF8FFFAFFFCFFFE0000",
		INIT_1B=>X"FFFE000100030005000600080009000A000A000A000900080006000500030001",
		INIT_1C=>X"00020000FFFEFFFCFFFAFFF8FFF7FFF6FFF5FFF5FFF5FFF6FFF7FFF9FFFAFFFC",
		INIT_1D=>X"FFFBFFFDFFFF00010004000500070009000A000A000A000A0009000800060004",
		INIT_1E=>X"000600040002FFFFFFFDFFFBFFF9FFF7FFF6FFF5FFF5FFF5FFF5FFF6FFF7FFF9",
		INIT_1F=>X"FFF8FFF9FFFBFFFE000000020004000600080009000A000B000B000A00090008",
		INIT_20=>X"00090007000500030001FFFFFFFCFFFAFFF8FFF6FFF5FFF4FFF4FFF4FFF5FFF6",
		INIT_21=>X"FFF5FFF6FFF8FFFAFFFCFFFE00010003000500070009000A000B000B000B000A",
		INIT_22=>X"000B000A00090007000500030000FFFEFFFBFFF9FFF7FFF6FFF4FFF4FFF4FFF4",
		INIT_23=>X"FFF3FFF3FFF5FFF6FFF8FFFAFFFDFFFF0002000400060008000A000B000C000C",
		INIT_24=>X"000C000C000C000B0009000700050002FFFFFFFDFFFAFFF8FFF6FFF5FFF3FFF3",
		INIT_25=>X"FFF2FFF2FFF2FFF3FFF4FFF6FFF8FFFBFFFD0000000300050008000A000B000C",
		INIT_26=>X"000C000D000D000D000C000B0009000700040001FFFEFFFCFFF9FFF7FFF5FFF3",
		INIT_27=>X"FFF4FFF2FFF1FFF1FFF2FFF3FFF4FFF6FFF9FFFBFFFE0001000400070009000B",
		INIT_28=>X"000A000C000D000E000E000E000D000B0009000600030000FFFDFFFAFFF8FFF5",
		INIT_29=>X"FFF6FFF4FFF2FFF1FFF0FFF0FFF1FFF2FFF4FFF6FFF9FFFCFFFF000200050008",
		INIT_2A=>X"0007000A000C000E000F000F000F000E000D000B000800060002FFFFFFFCFFF9",
		INIT_2B=>X"FFFBFFF7FFF5FFF2FFF0FFEFFFEFFFEFFFF0FFF2FFF4FFF7FFFAFFFD00000004",
		INIT_2C=>X"000200050009000B000E0010001100110010000F000E000B000800050002FFFE",
		INIT_2D=>X"0000FFFDFFF9FFF5FFF3FFF0FFEEFFEDFFEDFFEEFFEFFFF1FFF4FFF7FFFAFFFE",
		INIT_2E=>X"FFFBFFFF00030007000B000E001000120013001300120010000E000B00080004",
		INIT_2F=>X"00080003FFFFFFFBFFF7FFF3FFF0FFEEFFECFFEBFFEBFFECFFEEFFF1FFF4FFF7",
		INIT_30=>X"FFF4FFF8FFFC000100050009000D0010001300140015001500130011000F000B",
		INIT_31=>X"000F000B00070002FFFDFFF9FFF4FFF0FFEDFFEBFFE9FFE9FFE9FFEBFFEDFFF0",
		INIT_32=>X"FFEBFFEFFFF4FFF8FFFE00030008000C00100013001600170018001700150013",
		INIT_33=>X"001800150010000C00060001FFFBFFF6FFF1FFEDFFEAFFE7FFE6FFE6FFE7FFE8",
		INIT_34=>X"FFE3FFE6FFE9FFEEFFF3FFF9FFFF0005000B001000140018001A001B001B001A",
		INIT_35=>X"0020001E001B00170012000C0005FFFFFFF8FFF2FFEDFFE8FFE5FFE2FFE1FFE2",
		INIT_36=>X"FFDBFFDCFFDEFFE2FFE7FFEDFFF3FFFA00020009000F0015001A001D00200021",
		INIT_37=>X"00280028002700240020001A0013000C0004FFFCFFF4FFEDFFE7FFE2FFDEFFDC",
		INIT_38=>X"FFD4FFD2FFD2FFD3FFD7FFDCFFE3FFEBFFF3FFFC0005000E0015001C00220026",
		INIT_39=>X"002E0033003400340032002D0027001F0016000C0001FFF7FFEEFFE5FFDEFFD8",
		INIT_3A=>X"FFCEFFC7FFC3FFC1FFC2FFC5FFCBFFD3FFDDFFE8FFF3FFFF000B001600200028",
		INIT_3B=>X"0033003E0046004B004C004A0045003E00330027001A000CFFFDFFF0FFE3FFD7",
		INIT_3C=>X"FFCAFFB9FFACFFA3FF9EFF9DFFA1FFA8FFB3FFC0FFD0FFE1FFF3000500160026",
		INIT_3D=>X"003600520069007A0085008A00890082007600660052003C0024000CFFF4FFDE",
		INIT_3E=>X"FFC8FF8EFF5FFF3CFF24FF17FF15FF1DFF2DFF45FF62FF84FFA9FFCEFFF30016",
		INIT_3F=>X"04380430041903F303C00381033602E30289022A01C90168010900AE0059000C",
		INIT_40=>X"FFFFFFFDFFFBFFF9FFF8FFF8FFF8FFF9FFFAFFFCFFFE00000003000500060007",
		INIT_41=>X"FFF8FFF8FFFAFFFBFFFD00000002000400060007000700070007000500030001",
		INIT_42=>X"00010003000500070007000700070006000400020000FFFDFFFBFFF9FFF8FFF8",
		INIT_43=>X"00070006000500030000FFFEFFFCFFFAFFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF",
		INIT_44=>X"FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFAFFFCFFFE000100030005000600070008",
		INIT_45=>X"FFF8FFF9FFFBFFFD00000002000400060007000800070007000500030001FFFF",
		INIT_46=>X"0004000500070007000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF8",
		INIT_47=>X"0006000500030000FFFEFFFCFFFAFFF8FFF8FFF7FFF8FFF9FFFBFFFDFFFF0001",
		INIT_48=>X"FFFAFFF9FFF8FFF7FFF8FFF8FFFAFFFCFFFE0001000300050006000700080007",
		INIT_49=>X"FFF9FFFBFFFD00000002000400060007000800080007000500030001FFFFFFFD",
		INIT_4A=>X"000600070008000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF7FFF8",
		INIT_4B=>X"000500030000FFFEFFFCFFFAFFF8FFF7FFF7FFF8FFF9FFFBFFFDFFFF00010004",
		INIT_4C=>X"FFF9FFF8FFF7FFF7FFF8FFFAFFFCFFFE00010003000500070008000800070006",
		INIT_4D=>X"FFFBFFFD00000002000400060007000800080007000500030001FFFFFFFCFFFA",
		INIT_4E=>X"00070008000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF7FFF8FFF9",
		INIT_4F=>X"00030000FFFEFFFCFFFAFFF8FFF7FFF7FFF7FFF9FFFAFFFDFFFF000100040006",
		INIT_50=>X"FFF7FFF7FFF7FFF8FFFAFFFCFFFE000100030005000700080008000800070005",
		INIT_51=>X"FFFD00000002000500060008000800080007000600040001FFFFFFFCFFFAFFF8",
		INIT_52=>X"0008000800080006000400020000FFFDFFFBFFF9FFF7FFF7FFF7FFF8FFF9FFFB",
		INIT_53=>X"0000FFFEFFFBFFF9FFF8FFF7FFF6FFF7FFF8FFFAFFFCFFFF0002000400060008",
		INIT_54=>X"FFF6FFF7FFF8FFF9FFFCFFFE0001000300060007000800090008000700050003",
		INIT_55=>X"00000003000500070008000900090008000600040001FFFFFFFCFFFAFFF8FFF7",
		INIT_56=>X"00090008000700050002FFFFFFFDFFFAFFF8FFF7FFF6FFF6FFF7FFF9FFFBFFFD",
		INIT_57=>X"FFFEFFFBFFF9FFF7FFF6FFF6FFF7FFF8FFFAFFFCFFFF00020004000600080009",
		INIT_58=>X"FFF6FFF7FFF9FFFBFFFE00010004000600080009000900090007000600030000",
		INIT_59=>X"0003000500070009000900090008000600040001FFFFFFFCFFF9FFF7FFF6FFF6",
		INIT_5A=>X"0009000700050002FFFFFFFDFFFAFFF8FFF6FFF6FFF6FFF7FFF8FFFAFFFD0000",
		INIT_5B=>X"FFFBFFF8FFF6FFF5FFF5FFF6FFF7FFFAFFFCFFFF0002000500070009000A000A",
		INIT_5C=>X"FFF7FFF9FFFBFFFE0001000400070008000A000A00090008000600030000FFFD",
		INIT_5D=>X"00060008000A000A000A0009000700040001FFFEFFFBFFF9FFF7FFF5FFF5FFF5",
		INIT_5E=>X"000800050003FFFFFFFCFFF9FFF7FFF5FFF5FFF5FFF6FFF8FFFAFFFD00000003",
		INIT_5F=>X"FFF8FFF6FFF4FFF4FFF5FFF7FFF9FFFCFFFF000200050008000A000A000A000A",
		INIT_60=>X"FFF8FFFBFFFE0001000400070009000B000B000A0009000700040000FFFDFFFA",
		INIT_61=>X"0009000B000B000B000A000800050002FFFEFFFBFFF8FFF6FFF4FFF4FFF4FFF6",
		INIT_62=>X"00060003FFFFFFFCFFF9FFF6FFF4FFF3FFF4FFF5FFF7FFFAFFFD000000040007",
		INIT_63=>X"FFF4FFF3FFF3FFF4FFF6FFF8FFFCFFFF000300060009000B000C000C000B0009",
		INIT_64=>X"FFFAFFFE000200050008000B000C000C000C000A000700040001FFFDFFF9FFF7",
		INIT_65=>X"000C000D000D000B000900050002FFFEFFFAFFF7FFF5FFF3FFF2FFF3FFF5FFF7",
		INIT_66=>X"0003FFFFFFFBFFF8FFF5FFF3FFF2FFF2FFF3FFF6FFF9FFFD000000040008000A",
		INIT_67=>X"FFF1FFF1FFF2FFF4FFF7FFFBFFFF00030007000A000C000D000D000C000A0007",
		INIT_68=>X"FFFE00020006000A000C000E000E000D000B000800050001FFFCFFF8FFF5FFF3",
		INIT_69=>X"000F000F000D000A00060002FFFEFFF9FFF6FFF3FFF1FFF0FFF1FFF3FFF6FFF9",
		INIT_6A=>X"FFFFFFFAFFF6FFF3FFF1FFF0FFF0FFF1FFF4FFF8FFFC000100050009000C000E",
		INIT_6B=>X"FFEFFFF0FFF2FFF6FFFAFFFF00040008000C000F00100010000E000C00080004",
		INIT_6C=>X"00030007000C000F001100110010000E000A00060001FFFCFFF7FFF3FFF0FFEF",
		INIT_6D=>X"00120010000C00080003FFFDFFF8FFF4FFF0FFEEFFEDFFEEFFF0FFF4FFF8FFFD",
		INIT_6E=>X"FFF9FFF4FFF0FFEDFFECFFECFFEEFFF2FFF6FFFB00010006000B000F00110012",
		INIT_6F=>X"FFECFFEFFFF4FFF9FFFF0005000A000F0012001400130012000E000A0005FFFF",
		INIT_70=>X"0009000F00130015001500140011000D00070001FFFBFFF5FFF0FFEDFFEBFFEB",
		INIT_71=>X"0014000F000A0003FFFCFFF6FFF0FFECFFE9FFE9FFEAFFEDFFF1FFF7FFFD0003",
		INIT_72=>X"FFF1FFECFFE8FFE6FFE7FFEAFFEEFFF4FFFA00010008000E0013001600170017",
		INIT_73=>X"FFEAFFF0FFF7FFFF0007000E00140018001A001A00170013000D0006FFFFFFF7",
		INIT_74=>X"00140019001C001D001B0017001100090001FFF9FFF1FFEBFFE6FFE4FFE4FFE6",
		INIT_75=>X"0016000E0005FFFBFFF2FFEBFFE5FFE1FFE0FFE2FFE6FFECFFF4FFFC0005000D",
		INIT_76=>X"FFE3FFDEFFDCFFDCFFE0FFE7FFEFFFF80002000C0015001B001F00210020001C",
		INIT_77=>X"FFE9FFF4FFFF000B0015001D0023002600260022001C00130009FFFEFFF4FFEA",
		INIT_78=>X"0028002D002D002A0024001A000F0002FFF5FFEAFFE0FFD9FFD6FFD6FFD9FFE0",
		INIT_79=>X"00170008FFF8FFEAFFDDFFD4FFCEFFCDFFCFFFD6FFE0FFEDFFFA000800150020",
		INIT_7A=>X"FFC3FFBFFFC1FFC8FFD4FFE3FFF3000500160024002F003600380036002F0024",
		INIT_7B=>X"FFE8FFFF0016002A003A0045004A00480041003400240011FFFDFFE9FFD8FFCB",
		INIT_7C=>X"006A006A00610051003B00210005FFE9FFD1FFBDFFAFFFA8FFA9FFB1FFBFFFD2",
		INIT_7D=>X"0017FFE9FFBFFF9DFF85FF78FF76FF80FF94FFB0FFD0FFF300160035004E0060",
		INIT_7E=>X"FEBAFED4FF02FF3FFF86FFCF00160055008700AB00BE00C100B3009900730047",
		INIT_7F=>X"05E805D20594053004AB040B0358029C01DD0126007DFFE9FF70FF14FED8FEBB",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_08,
		DOPADOP=>dopadop_08,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_09: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"00FFFFFC00000FFFFF000003FFFFF000003FFFFF000003FFFFC00000FFFFFC00",
		INITP_01=>X"0FFFFFC00000FFFFF000003FFFFF000003FFFFF000003FFFFC00000FFFFFC000",
		INITP_02=>X"FFFFFC00003FFFFF000003FFFFF000003FFFFF000003FFFFC00000FFFFFC0000",
		INITP_03=>X"FFFFC00003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000",
		INITP_04=>X"FFFC00003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000F",
		INITP_05=>X"FFC00003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000FF",
		INITP_06=>X"FC00003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000FFF",
		INITP_07=>X"000003FFFFF000003FFFFF000003FFFFF00000FFFFFC00000FFFFFC00000FFFF",
		INITP_08=>X"0FFFF0003FFFC0003FFF0000FFFF0003FFFC0003FFF0000FFFF0003FFFC0003F",
		INITP_09=>X"0003FFFC0003FFF0000FFFF0003FFFC0003FFF0000FFFF0003FFFC0003FFF000",
		INITP_0A=>X"FFC000FFFF0000FFFC0003FFFC0003FFF0000FFFF0003FFFC0003FFF0000FFFF",
		INITP_0B=>X"0FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003F",
		INITP_0C=>X"0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC00",
		INITP_0D=>X"FFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF",
		INITP_0E=>X"03FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000F",
		INITP_0F=>X"0000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC00",
		INIT_00=>X"FFFFFFFDFFFBFFF9FFF8FFF8FFF8FFF9FFFAFFFCFFFE00000003000500060007",
		INIT_01=>X"FFF8FFF8FFFAFFFBFFFD00000002000400060007000700070007000500030001",
		INIT_02=>X"00010003000500070007000700070006000400020000FFFDFFFBFFF9FFF8FFF8",
		INIT_03=>X"00070006000500030000FFFEFFFCFFFAFFF9FFF8FFF7FFF8FFF9FFFBFFFDFFFF",
		INIT_04=>X"FFFDFFFBFFF9FFF8FFF7FFF8FFF9FFFAFFFCFFFE000100030005000600070008",
		INIT_05=>X"FFF8FFF9FFFBFFFD00000002000400060007000800070007000500030001FFFF",
		INIT_06=>X"0004000500070007000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF8",
		INIT_07=>X"0006000500030000FFFEFFFCFFFAFFF8FFF8FFF7FFF8FFF9FFFBFFFDFFFF0001",
		INIT_08=>X"FFFAFFF9FFF8FFF7FFF8FFF8FFFAFFFCFFFE0001000300050006000700080007",
		INIT_09=>X"FFF9FFFBFFFD00000002000400060007000800080007000500030001FFFFFFFD",
		INIT_0A=>X"000600070008000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF7FFF8",
		INIT_0B=>X"000500030000FFFEFFFCFFFAFFF8FFF7FFF7FFF8FFF9FFFBFFFDFFFF00010004",
		INIT_0C=>X"FFF9FFF8FFF7FFF7FFF8FFFAFFFCFFFE00010003000500070008000800070006",
		INIT_0D=>X"FFFBFFFD00000002000400060007000800080007000500030001FFFFFFFCFFFA",
		INIT_0E=>X"00070008000800070006000400020000FFFDFFFBFFF9FFF8FFF7FFF7FFF8FFF9",
		INIT_0F=>X"00030000FFFEFFFCFFFAFFF8FFF7FFF7FFF7FFF9FFFAFFFDFFFF000100040006",
		INIT_10=>X"FFF7FFF7FFF7FFF8FFFAFFFCFFFE000100030005000700080008000800070005",
		INIT_11=>X"FFFD00000002000500060008000800080007000600040001FFFFFFFCFFFAFFF8",
		INIT_12=>X"0008000800080006000400020000FFFDFFFBFFF9FFF7FFF7FFF7FFF8FFF9FFFB",
		INIT_13=>X"0000FFFEFFFBFFF9FFF8FFF7FFF6FFF7FFF8FFFAFFFCFFFF0002000400060008",
		INIT_14=>X"FFF6FFF7FFF8FFF9FFFCFFFE0001000300060007000800090008000700050003",
		INIT_15=>X"00000003000500070008000900090008000600040001FFFFFFFCFFFAFFF8FFF7",
		INIT_16=>X"00090008000700050002FFFFFFFDFFFAFFF8FFF7FFF6FFF6FFF7FFF9FFFBFFFD",
		INIT_17=>X"FFFEFFFBFFF9FFF7FFF6FFF6FFF7FFF8FFFAFFFCFFFF00020004000600080009",
		INIT_18=>X"FFF6FFF7FFF9FFFBFFFE00010004000600080009000900090007000600030000",
		INIT_19=>X"0003000500070009000900090008000600040001FFFFFFFCFFF9FFF7FFF6FFF6",
		INIT_1A=>X"0009000700050002FFFFFFFDFFFAFFF8FFF6FFF6FFF6FFF7FFF8FFFAFFFD0000",
		INIT_1B=>X"FFFBFFF8FFF6FFF5FFF5FFF6FFF7FFFAFFFCFFFF0002000500070009000A000A",
		INIT_1C=>X"FFF7FFF9FFFBFFFE0001000400070008000A000A00090008000600030000FFFD",
		INIT_1D=>X"00060008000A000A000A0009000700040001FFFEFFFBFFF9FFF7FFF5FFF5FFF5",
		INIT_1E=>X"000800050003FFFFFFFCFFF9FFF7FFF5FFF5FFF5FFF6FFF8FFFAFFFD00000003",
		INIT_1F=>X"FFF8FFF6FFF4FFF4FFF5FFF7FFF9FFFCFFFF000200050008000A000A000A000A",
		INIT_20=>X"FFF8FFFBFFFE0001000400070009000B000B000A0009000700040000FFFDFFFA",
		INIT_21=>X"0009000B000B000B000A000800050002FFFEFFFBFFF8FFF6FFF4FFF4FFF4FFF6",
		INIT_22=>X"00060003FFFFFFFCFFF9FFF6FFF4FFF3FFF4FFF5FFF7FFFAFFFD000000040007",
		INIT_23=>X"FFF4FFF3FFF3FFF4FFF6FFF8FFFCFFFF000300060009000B000C000C000B0009",
		INIT_24=>X"FFFAFFFE000200050008000B000C000C000C000A000700040001FFFDFFF9FFF7",
		INIT_25=>X"000C000D000D000B000900050002FFFEFFFAFFF7FFF5FFF3FFF2FFF3FFF5FFF7",
		INIT_26=>X"0003FFFFFFFBFFF8FFF5FFF3FFF2FFF2FFF3FFF6FFF9FFFD000000040008000A",
		INIT_27=>X"FFF1FFF1FFF2FFF4FFF7FFFBFFFF00030007000A000C000D000D000C000A0007",
		INIT_28=>X"FFFE00020006000A000C000E000E000D000B000800050001FFFCFFF8FFF5FFF3",
		INIT_29=>X"000F000F000D000A00060002FFFEFFF9FFF6FFF3FFF1FFF0FFF1FFF3FFF6FFF9",
		INIT_2A=>X"FFFFFFFAFFF6FFF3FFF1FFF0FFF0FFF1FFF4FFF8FFFC000100050009000C000E",
		INIT_2B=>X"FFEFFFF0FFF2FFF6FFFAFFFF00040008000C000F00100010000E000C00080004",
		INIT_2C=>X"00030007000C000F001100110010000E000A00060001FFFCFFF7FFF3FFF0FFEF",
		INIT_2D=>X"00120010000C00080003FFFDFFF8FFF4FFF0FFEEFFEDFFEEFFF0FFF4FFF8FFFD",
		INIT_2E=>X"FFF9FFF4FFF0FFEDFFECFFECFFEEFFF2FFF6FFFB00010006000B000F00110012",
		INIT_2F=>X"FFECFFEFFFF4FFF9FFFF0005000A000F0012001400130012000E000A0005FFFF",
		INIT_30=>X"0009000F00130015001500140011000D00070001FFFBFFF5FFF0FFEDFFEBFFEB",
		INIT_31=>X"0014000F000A0003FFFCFFF6FFF0FFECFFE9FFE9FFEAFFEDFFF1FFF7FFFD0003",
		INIT_32=>X"FFF1FFECFFE8FFE6FFE7FFEAFFEEFFF4FFFA00010008000E0013001600170017",
		INIT_33=>X"FFEAFFF0FFF7FFFF0007000E00140018001A001A00170013000D0006FFFFFFF7",
		INIT_34=>X"00140019001C001D001B0017001100090001FFF9FFF1FFEBFFE6FFE4FFE4FFE6",
		INIT_35=>X"0016000E0005FFFBFFF2FFEBFFE5FFE1FFE0FFE2FFE6FFECFFF4FFFC0005000D",
		INIT_36=>X"FFE3FFDEFFDCFFDCFFE0FFE7FFEFFFF80002000C0015001B001F00210020001C",
		INIT_37=>X"FFE9FFF4FFFF000B0015001D0023002600260022001C00130009FFFEFFF4FFEA",
		INIT_38=>X"0028002D002D002A0024001A000F0002FFF5FFEAFFE0FFD9FFD6FFD6FFD9FFE0",
		INIT_39=>X"00170008FFF8FFEAFFDDFFD4FFCEFFCDFFCFFFD6FFE0FFEDFFFA000800150020",
		INIT_3A=>X"FFC3FFBFFFC1FFC8FFD4FFE3FFF3000500160024002F003600380036002F0024",
		INIT_3B=>X"FFE8FFFF0016002A003A0045004A00480041003400240011FFFDFFE9FFD8FFCB",
		INIT_3C=>X"006A006A00610051003B00210005FFE9FFD1FFBDFFAFFFA8FFA9FFB1FFBFFFD2",
		INIT_3D=>X"0017FFE9FFBFFF9DFF85FF78FF76FF80FF94FFB0FFD0FFF300160035004E0060",
		INIT_3E=>X"FEBAFED4FF02FF3FFF86FFCF00160055008700AB00BE00C100B3009900730047",
		INIT_3F=>X"05E805D20594053004AB040B0358029C01DD0126007DFFE9FF70FF14FED8FEBB",
		INIT_40=>X"FFF8FFF8FFF9FFFBFFFE00010004000600070007000600030000FFFDFFFAFFF8",
		INIT_41=>X"FFF9FFF8FFF8FFF9FFFCFFFF0002000500070008000700050002FFFFFFFCFFF9",
		INIT_42=>X"FFFAFFF8FFF7FFF8FFFAFFFD00000003000600070007000600040001FFFEFFFB",
		INIT_43=>X"FFFCFFF9FFF8FFF8FFF9FFFBFFFE00010004000600070007000600030000FFFD",
		INIT_44=>X"FFFEFFFBFFF9FFF8FFF8FFF9FFFCFFFF0002000500070008000700050002FFFF",
		INIT_45=>X"0000FFFDFFFAFFF8FFF7FFF8FFFAFFFD00000003000600070007000600040001",
		INIT_46=>X"0002FFFFFFFCFFF9FFF8FFF7FFF9FFFBFFFE0001000400070008000700060003",
		INIT_47=>X"00040001FFFEFFFBFFF8FFF7FFF8FFF9FFFCFFFF000200050007000800070005",
		INIT_48=>X"000600030000FFFDFFFAFFF8FFF7FFF8FFFAFFFD000000030006000700080006",
		INIT_49=>X"000700050002FFFFFFFBFFF9FFF8FFF7FFF9FFFBFFFE00010004000700080007",
		INIT_4A=>X"0008000600040001FFFEFFFAFFF8FFF7FFF8FFF9FFFCFFFF0003000500070008",
		INIT_4B=>X"00080007000600030000FFFCFFFAFFF8FFF7FFF8FFFAFFFD0000000400060008",
		INIT_4C=>X"00070008000700050002FFFFFFFBFFF9FFF7FFF7FFF9FFFBFFFE000200050007",
		INIT_4D=>X"000600080008000700040001FFFDFFFAFFF8FFF7FFF7FFF9FFFCFFFF00030006",
		INIT_4E=>X"0005000700080008000600030000FFFCFFF9FFF8FFF7FFF8FFFAFFFD00000004",
		INIT_4F=>X"0003000600080008000700050002FFFEFFFBFFF9FFF7FFF7FFF8FFFBFFFE0002",
		INIT_50=>X"00010004000700080008000700040001FFFDFFFAFFF8FFF7FFF7FFF9FFFCFFFF",
		INIT_51=>X"FFFE00020005000700080008000600030000FFFCFFF9FFF7FFF7FFF8FFFAFFFD",
		INIT_52=>X"FFFCFFFF0003000600080008000700050002FFFEFFFBFFF8FFF7FFF7FFF8FFFB",
		INIT_53=>X"FFFAFFFD00010004000700080008000700040001FFFDFFFAFFF8FFF7FFF7FFF9",
		INIT_54=>X"FFF8FFFBFFFE00020005000800090008000600030000FFFCFFF9FFF7FFF6FFF7",
		INIT_55=>X"FFF7FFF9FFFC00000003000600080009000800050002FFFEFFFBFFF8FFF6FFF6",
		INIT_56=>X"FFF6FFF7FFFAFFFD00010004000700090009000700040001FFFDFFFAFFF7FFF6",
		INIT_57=>X"FFF6FFF6FFF8FFFBFFFE0002000600080009000800060003FFFFFFFCFFF9FFF7",
		INIT_58=>X"FFF7FFF6FFF6FFF8FFFC00000003000700090009000800060002FFFEFFFAFFF8",
		INIT_59=>X"FFF8FFF6FFF6FFF7FFF9FFFD00010005000800090009000700050001FFFDFFF9",
		INIT_5A=>X"FFFAFFF7FFF6FFF6FFF7FFFAFFFE000200060008000A000900070003FFFFFFFB",
		INIT_5B=>X"FFFCFFF9FFF6FFF5FFF6FFF8FFFC0000000400070009000A000800060002FFFE",
		INIT_5C=>X"FFFFFFFBFFF8FFF6FFF5FFF6FFF9FFFD000100050008000A000A000800050001",
		INIT_5D=>X"0002FFFEFFFAFFF7FFF5FFF5FFF7FFFAFFFE000300060009000A000900070003",
		INIT_5E=>X"00050001FFFCFFF8FFF6FFF5FFF5FFF8FFFB000000040008000A000A00090006",
		INIT_5F=>X"00080004FFFFFFFBFFF7FFF5FFF4FFF6FFF9FFFD000100060009000A000A0008",
		INIT_60=>X"000A00060002FFFEFFF9FFF6FFF4FFF4FFF6FFFAFFFE00030007000A000B000A",
		INIT_61=>X"000B000900050001FFFCFFF8FFF5FFF4FFF5FFF7FFFB000000050008000B000B",
		INIT_62=>X"000C000B00080004FFFFFFFAFFF6FFF4FFF3FFF5FFF8FFFD00020006000A000B",
		INIT_63=>X"000C000C000A00070002FFFDFFF9FFF5FFF3FFF3FFF6FFFAFFFE00030008000B",
		INIT_64=>X"000A000C000C000A00060001FFFBFFF7FFF4FFF3FFF4FFF7FFFB000000050009",
		INIT_65=>X"0009000C000D000C00090004FFFFFFFAFFF5FFF3FFF2FFF4FFF8FFFD00020007",
		INIT_66=>X"0006000A000D000D000B00080002FFFDFFF8FFF4FFF2FFF2FFF5FFF9FFFE0004",
		INIT_67=>X"00020008000C000E000D000B00060001FFFBFFF6FFF3FFF1FFF3FFF6FFFB0000",
		INIT_68=>X"FFFE0004000A000D000E000D000A0005FFFFFFF9FFF4FFF2FFF1FFF3FFF7FFFC",
		INIT_69=>X"FFFA00010007000B000E000F000D00080003FFFCFFF7FFF3FFF1FFF1FFF4FFF9",
		INIT_6A=>X"FFF6FFFC00030009000D000F000F000C00070001FFFAFFF5FFF1FFF0FFF1FFF5",
		INIT_6B=>X"FFF2FFF8FFFE0005000B000F0010000F000B0005FFFEFFF8FFF3FFF0FFEFFFF2",
		INIT_6C=>X"FFEFFFF3FFFA00010008000D00100011000E00090003FFFCFFF6FFF1FFEFFFEF",
		INIT_6D=>X"FFEDFFF0FFF5FFFC0003000A000F00120011000E00080001FFF9FFF3FFEFFFEE",
		INIT_6E=>X"FFECFFEDFFF0FFF7FFFE0006000D001100130011000C0006FFFEFFF7FFF1FFED",
		INIT_6F=>X"FFECFFEBFFEDFFF2FFF9000100090010001300130011000B0003FFFBFFF4FFEE",
		INIT_70=>X"FFEEFFEAFFEAFFEDFFF3FFFB0004000C001200150014001000090001FFF8FFF1",
		INIT_71=>X"FFF1FFEBFFE8FFE9FFEEFFF5FFFE00080010001500160014000F0007FFFEFFF5",
		INIT_72=>X"FFF6FFEEFFE8FFE6FFE9FFEFFFF80002000B0013001700170014000D0004FFFA",
		INIT_73=>X"FFFDFFF2FFEAFFE5FFE5FFE9FFF1FFFB0006000F0016001900180013000B0001",
		INIT_74=>X"0005FFF8FFEEFFE6FFE2FFE4FFEAFFF3FFFE000A0014001A001C001900120008",
		INIT_75=>X"000E0001FFF4FFE9FFE2FFE0FFE3FFEBFFF60003000F0018001D001E00190010",
		INIT_76=>X"0017000AFFFCFFEEFFE3FFDDFFDDFFE2FFEDFFFA00080014001D0021001F0018",
		INIT_77=>X"002200160006FFF6FFE7FFDDFFD8FFDAFFE3FFEFFFFE000E001A002200240021",
		INIT_78=>X"002C002200130001FFEEFFDFFFD6FFD3FFD8FFE3FFF300040015002100280028",
		INIT_79=>X"003600300022000FFFF9FFE5FFD6FFCEFFCEFFD6FFE5FFF8000C001D0029002F",
		INIT_7A=>X"003F003F003400210009FFF0FFDAFFCBFFC4FFC8FFD4FFE8FFFE001500270033",
		INIT_7B=>X"00470050004A0039001F0001FFE3FFCAFFBBFFB8FFC0FFD3FFEC000800210035",
		INIT_7C=>X"004E00640068005B0040001BFFF3FFCFFFB4FFA6FFA7FFB7FFD1FFF300150033",
		INIT_7D=>X"00530080009600920077004A0013FFDCFFAEFF8FFF84FF8DFFA8FFD0FFFE002B",
		INIT_7E=>X"005600C00100011100F600B6005F0001FFAAFF68FF43FF3FFF5AFF8DFFD00015",
		INIT_7F=>X"0858081C077106650514039E022500CAFFA8FED3FE56FE2FFE56FEB7FF3DFFCF",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_09,
		DOPADOP=>dopadop_09,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_10: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"0FFFF0003FFFC0003FFF0000FFFF0003FFFC0003FFF0000FFFF0003FFFC0003F",
		INITP_01=>X"0003FFFC0003FFF0000FFFF0003FFFC0003FFF0000FFFF0003FFFC0003FFF000",
		INITP_02=>X"FFC000FFFF0000FFFC0003FFFC0003FFF0000FFFF0003FFFC0003FFF0000FFFF",
		INITP_03=>X"0FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003F",
		INITP_04=>X"0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC00",
		INITP_05=>X"FFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF",
		INITP_06=>X"03FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000F",
		INITP_07=>X"0000FFFF0000FFFC0003FFFC000FFFF0000FFFC0003FFFC000FFFF0000FFFC00",
		INITP_08=>X"000FFC003FF003FFC00FFF003FFC00FFF003FFC00FFF003FF000FFC003FF000F",
		INITP_09=>X"03FF003FFC00FFF003FFC00FFF003FFC00FFF003FF000FFC003FF000FFC003FF",
		INITP_0A=>X"FFC00FFF003FFC00FFF003FFC00FFF003FF000FFC003FF000FFC003FF000FFC0",
		INITP_0B=>X"F003FFC00FFF003FFC00FFF003FF000FFC003FF000FFC003FF000FFC003FF003",
		INITP_0C=>X"00FFF003FFC00FFF003FF000FFC003FF000FFC003FF000FFC003FF003FFC00FF",
		INITP_0D=>X"3FFC00FFF003FF000FFC003FF000FFC003FF000FFC003FF003FFC00FFF003FFC",
		INITP_0E=>X"FF003FF000FFC003FF000FFC003FF000FFC003FF003FFC00FFF003FFC00FFF00",
		INITP_0F=>X"000FFC003FF000FFC003FF000FFC003FF003FFC00FFF003FFC00FFF003FFC00F",
		INIT_00=>X"FFF8FFF8FFF9FFFBFFFE00010004000600070007000600030000FFFDFFFAFFF8",
		INIT_01=>X"FFF9FFF8FFF8FFF9FFFCFFFF0002000500070008000700050002FFFFFFFCFFF9",
		INIT_02=>X"FFFAFFF8FFF7FFF8FFFAFFFD00000003000600070007000600040001FFFEFFFB",
		INIT_03=>X"FFFCFFF9FFF8FFF8FFF9FFFBFFFE00010004000600070007000600030000FFFD",
		INIT_04=>X"FFFEFFFBFFF9FFF8FFF8FFF9FFFCFFFF0002000500070008000700050002FFFF",
		INIT_05=>X"0000FFFDFFFAFFF8FFF7FFF8FFFAFFFD00000003000600070007000600040001",
		INIT_06=>X"0002FFFFFFFCFFF9FFF8FFF7FFF9FFFBFFFE0001000400070008000700060003",
		INIT_07=>X"00040001FFFEFFFBFFF8FFF7FFF8FFF9FFFCFFFF000200050007000800070005",
		INIT_08=>X"000600030000FFFDFFFAFFF8FFF7FFF8FFFAFFFD000000030006000700080006",
		INIT_09=>X"000700050002FFFFFFFBFFF9FFF8FFF7FFF9FFFBFFFE00010004000700080007",
		INIT_0A=>X"0008000600040001FFFEFFFAFFF8FFF7FFF8FFF9FFFCFFFF0003000500070008",
		INIT_0B=>X"00080007000600030000FFFCFFFAFFF8FFF7FFF8FFFAFFFD0000000400060008",
		INIT_0C=>X"00070008000700050002FFFFFFFBFFF9FFF7FFF7FFF9FFFBFFFE000200050007",
		INIT_0D=>X"000600080008000700040001FFFDFFFAFFF8FFF7FFF7FFF9FFFCFFFF00030006",
		INIT_0E=>X"0005000700080008000600030000FFFCFFF9FFF8FFF7FFF8FFFAFFFD00000004",
		INIT_0F=>X"0003000600080008000700050002FFFEFFFBFFF9FFF7FFF7FFF8FFFBFFFE0002",
		INIT_10=>X"00010004000700080008000700040001FFFDFFFAFFF8FFF7FFF7FFF9FFFCFFFF",
		INIT_11=>X"FFFE00020005000700080008000600030000FFFCFFF9FFF7FFF7FFF8FFFAFFFD",
		INIT_12=>X"FFFCFFFF0003000600080008000700050002FFFEFFFBFFF8FFF7FFF7FFF8FFFB",
		INIT_13=>X"FFFAFFFD00010004000700080008000700040001FFFDFFFAFFF8FFF7FFF7FFF9",
		INIT_14=>X"FFF8FFFBFFFE00020005000800090008000600030000FFFCFFF9FFF7FFF6FFF7",
		INIT_15=>X"FFF7FFF9FFFC00000003000600080009000800050002FFFEFFFBFFF8FFF6FFF6",
		INIT_16=>X"FFF6FFF7FFFAFFFD00010004000700090009000700040001FFFDFFFAFFF7FFF6",
		INIT_17=>X"FFF6FFF6FFF8FFFBFFFE0002000600080009000800060003FFFFFFFCFFF9FFF7",
		INIT_18=>X"FFF7FFF6FFF6FFF8FFFC00000003000700090009000800060002FFFEFFFAFFF8",
		INIT_19=>X"FFF8FFF6FFF6FFF7FFF9FFFD00010005000800090009000700050001FFFDFFF9",
		INIT_1A=>X"FFFAFFF7FFF6FFF6FFF7FFFAFFFE000200060008000A000900070003FFFFFFFB",
		INIT_1B=>X"FFFCFFF9FFF6FFF5FFF6FFF8FFFC0000000400070009000A000800060002FFFE",
		INIT_1C=>X"FFFFFFFBFFF8FFF6FFF5FFF6FFF9FFFD000100050008000A000A000800050001",
		INIT_1D=>X"0002FFFEFFFAFFF7FFF5FFF5FFF7FFFAFFFE000300060009000A000900070003",
		INIT_1E=>X"00050001FFFCFFF8FFF6FFF5FFF5FFF8FFFB000000040008000A000A00090006",
		INIT_1F=>X"00080004FFFFFFFBFFF7FFF5FFF4FFF6FFF9FFFD000100060009000A000A0008",
		INIT_20=>X"000A00060002FFFEFFF9FFF6FFF4FFF4FFF6FFFAFFFE00030007000A000B000A",
		INIT_21=>X"000B000900050001FFFCFFF8FFF5FFF4FFF5FFF7FFFB000000050008000B000B",
		INIT_22=>X"000C000B00080004FFFFFFFAFFF6FFF4FFF3FFF5FFF8FFFD00020006000A000B",
		INIT_23=>X"000C000C000A00070002FFFDFFF9FFF5FFF3FFF3FFF6FFFAFFFE00030008000B",
		INIT_24=>X"000A000C000C000A00060001FFFBFFF7FFF4FFF3FFF4FFF7FFFB000000050009",
		INIT_25=>X"0009000C000D000C00090004FFFFFFFAFFF5FFF3FFF2FFF4FFF8FFFD00020007",
		INIT_26=>X"0006000A000D000D000B00080002FFFDFFF8FFF4FFF2FFF2FFF5FFF9FFFE0004",
		INIT_27=>X"00020008000C000E000D000B00060001FFFBFFF6FFF3FFF1FFF3FFF6FFFB0000",
		INIT_28=>X"FFFE0004000A000D000E000D000A0005FFFFFFF9FFF4FFF2FFF1FFF3FFF7FFFC",
		INIT_29=>X"FFFA00010007000B000E000F000D00080003FFFCFFF7FFF3FFF1FFF1FFF4FFF9",
		INIT_2A=>X"FFF6FFFC00030009000D000F000F000C00070001FFFAFFF5FFF1FFF0FFF1FFF5",
		INIT_2B=>X"FFF2FFF8FFFE0005000B000F0010000F000B0005FFFEFFF8FFF3FFF0FFEFFFF2",
		INIT_2C=>X"FFEFFFF3FFFA00010008000D00100011000E00090003FFFCFFF6FFF1FFEFFFEF",
		INIT_2D=>X"FFEDFFF0FFF5FFFC0003000A000F00120011000E00080001FFF9FFF3FFEFFFEE",
		INIT_2E=>X"FFECFFEDFFF0FFF7FFFE0006000D001100130011000C0006FFFEFFF7FFF1FFED",
		INIT_2F=>X"FFECFFEBFFEDFFF2FFF9000100090010001300130011000B0003FFFBFFF4FFEE",
		INIT_30=>X"FFEEFFEAFFEAFFEDFFF3FFFB0004000C001200150014001000090001FFF8FFF1",
		INIT_31=>X"FFF1FFEBFFE8FFE9FFEEFFF5FFFE00080010001500160014000F0007FFFEFFF5",
		INIT_32=>X"FFF6FFEEFFE8FFE6FFE9FFEFFFF80002000B0013001700170014000D0004FFFA",
		INIT_33=>X"FFFDFFF2FFEAFFE5FFE5FFE9FFF1FFFB0006000F0016001900180013000B0001",
		INIT_34=>X"0005FFF8FFEEFFE6FFE2FFE4FFEAFFF3FFFE000A0014001A001C001900120008",
		INIT_35=>X"000E0001FFF4FFE9FFE2FFE0FFE3FFEBFFF60003000F0018001D001E00190010",
		INIT_36=>X"0017000AFFFCFFEEFFE3FFDDFFDDFFE2FFEDFFFA00080014001D0021001F0018",
		INIT_37=>X"002200160006FFF6FFE7FFDDFFD8FFDAFFE3FFEFFFFE000E001A002200240021",
		INIT_38=>X"002C002200130001FFEEFFDFFFD6FFD3FFD8FFE3FFF300040015002100280028",
		INIT_39=>X"003600300022000FFFF9FFE5FFD6FFCEFFCEFFD6FFE5FFF8000C001D0029002F",
		INIT_3A=>X"003F003F003400210009FFF0FFDAFFCBFFC4FFC8FFD4FFE8FFFE001500270033",
		INIT_3B=>X"00470050004A0039001F0001FFE3FFCAFFBBFFB8FFC0FFD3FFEC000800210035",
		INIT_3C=>X"004E00640068005B0040001BFFF3FFCFFFB4FFA6FFA7FFB7FFD1FFF300150033",
		INIT_3D=>X"00530080009600920077004A0013FFDCFFAEFF8FFF84FF8DFFA8FFD0FFFE002B",
		INIT_3E=>X"005600C00100011100F600B6005F0001FFAAFF68FF43FF3FFF5AFF8DFFD00015",
		INIT_3F=>X"0858081C077106650514039E022500CAFFA8FED3FE56FE2FFE56FEB7FF3DFFCF",
		INIT_40=>X"000700050001FFFDFFF9FFF8FFF9FFFC000000050007000700050001FFFCFFF9",
		INIT_41=>X"FFF8FFFB000000040007000700050001FFFDFFF9FFF8FFF8FFFC000000040007",
		INIT_42=>X"00060002FFFEFFFAFFF8FFF8FFFBFFFF00040007000700060002FFFDFFF9FFF8",
		INIT_43=>X"FFFAFFFF00030006000800060002FFFEFFFAFFF8FFF8FFFBFFFF000300070007",
		INIT_44=>X"0003FFFFFFFAFFF8FFF8FFFAFFFE00030006000800060003FFFEFFFAFFF8FFF8",
		INIT_45=>X"FFFE00020006000800070003FFFFFFFBFFF8FFF8FFFAFFFE0002000600080006",
		INIT_46=>X"0000FFFBFFF8FFF7FFF9FFFD00020006000800070004FFFFFFFBFFF8FFF8FFFA",
		INIT_47=>X"000100050007000700040000FFFCFFF8FFF7FFF9FFFD00010005000700070004",
		INIT_48=>X"FFFCFFF9FFF7FFF9FFFC000100050007000700050000FFFCFFF8FFF7FFF9FFFC",
		INIT_49=>X"00040007000800050001FFFDFFF9FFF7FFF8FFFC000000050007000700050001",
		INIT_4A=>X"FFF9FFF7FFF8FFFB000000040007000800060002FFFDFFF9FFF7FFF8FFFB0000",
		INIT_4B=>X"0007000800060002FFFEFFF9FFF7FFF8FFFBFFFF00040007000800060002FFFD",
		INIT_4C=>X"FFF7FFF7FFFAFFFF00030007000800060003FFFEFFFAFFF7FFF8FFFAFFFF0004",
		INIT_4D=>X"000800070003FFFFFFFAFFF7FFF7FFFAFFFE00030007000800070003FFFEFFFA",
		INIT_4E=>X"FFF7FFF9FFFD00020006000800070004FFFFFFFAFFF8FFF7FFFAFFFE00030006",
		INIT_4F=>X"000800040000FFFBFFF8FFF7FFF9FFFD00020006000800070004FFFFFFFBFFF8",
		INIT_50=>X"FFF8FFFC000100060008000800050000FFFBFFF8FFF7FFF9FFFD000200060008",
		INIT_51=>X"00050001FFFCFFF8FFF7FFF8FFFC000100050008000800050001FFFCFFF8FFF7",
		INIT_52=>X"FFFB000000050008000800060001FFFCFFF8FFF7FFF8FFFB0000000500080008",
		INIT_53=>X"0002FFFDFFF9FFF7FFF7FFFB000000050008000800060002FFFDFFF8FFF7FFF8",
		INIT_54=>X"FFFF00040008000900070003FFFDFFF9FFF7FFF7FFFAFFFF0004000800090006",
		INIT_55=>X"FFFEFFF9FFF7FFF7FFFAFFFE00040007000900070003FFFEFFF9FFF7FFF7FFFA",
		INIT_56=>X"00030007000900080004FFFFFFFAFFF7FFF6FFF9FFFE00030007000900070003",
		INIT_57=>X"FFFAFFF7FFF6FFF8FFFD00030007000900080004FFFFFFFAFFF7FFF6FFF9FFFE",
		INIT_58=>X"00070009000900050000FFFAFFF7FFF6FFF8FFFD00020007000900080005FFFF",
		INIT_59=>X"FFF7FFF6FFF7FFFC000100060009000900050000FFFBFFF7FFF6FFF8FFFC0002",
		INIT_5A=>X"0009000900060001FFFBFFF7FFF5FFF7FFFB000100060009000900060001FFFB",
		INIT_5B=>X"FFF5FFF6FFFA000000060009000A00070002FFFCFFF7FFF5FFF7FFFB00010006",
		INIT_5C=>X"000A00080003FFFDFFF8FFF5FFF6FFFA000000050009000A00070002FFFCFFF7",
		INIT_5D=>X"FFF5FFF9FFFF00050009000A00080003FFFDFFF8FFF5FFF6FFF9FFFF00050009",
		INIT_5E=>X"00090004FFFEFFF8FFF5FFF5FFF8FFFE00040009000A00080004FFFDFFF8FFF5",
		INIT_5F=>X"FFF8FFFD00040009000B00090005FFFEFFF9FFF5FFF5FFF8FFFE00040009000B",
		INIT_60=>X"0006FFFFFFF9FFF5FFF4FFF7FFFD00030008000B000A0005FFFFFFF9FFF5FFF4",
		INIT_61=>X"FFFB00020008000B000A00060000FFF9FFF5FFF4FFF7FFFC00030008000B000A",
		INIT_62=>X"0001FFFAFFF5FFF3FFF6FFFB00020008000B000B00070000FFFAFFF5FFF4FFF6",
		INIT_63=>X"00010007000B000C00080002FFFBFFF5FFF3FFF5FFFA00010008000B000B0007",
		INIT_64=>X"FFFBFFF5FFF3FFF4FFF900000007000B000C00090002FFFBFFF5FFF3FFF5FFFA",
		INIT_65=>X"0006000C000D000A0003FFFCFFF6FFF2FFF3FFF800000007000C000C00090003",
		INIT_66=>X"FFF6FFF2FFF2FFF7FFFE0006000C000D000A0004FFFCFFF6FFF2FFF3FFF8FFFF",
		INIT_67=>X"000B000E000C0006FFFDFFF6FFF2FFF2FFF6FFFE0006000C000E000B0005FFFD",
		INIT_68=>X"FFF2FFF1FFF5FFFC0005000B000E000C0006FFFEFFF6FFF2FFF1FFF6FFFD0005",
		INIT_69=>X"000F000E0008FFFFFFF7FFF1FFF0FFF4FFFC0004000B000F000D0007FFFFFFF7",
		INIT_6A=>X"FFEFFFF3FFFA0003000B000F000E00090000FFF7FFF1FFF0FFF3FFFB0004000B",
		INIT_6B=>X"0010000A0002FFF8FFF1FFEFFFF2FFF90003000B0010000F000A0001FFF8FFF1",
		INIT_6C=>X"FFF0FFF70001000A00100010000B0002FFF9FFF1FFEEFFF1FFF80002000B0010",
		INIT_6D=>X"000D0004FFFAFFF1FFEDFFEFFFF60000000A00100011000C0003FFF9FFF1FFEE",
		INIT_6E=>X"FFF4FFFF000A00110013000E0005FFFAFFF1FFEDFFEEFFF50000000A00110012",
		INIT_6F=>X"0008FFFCFFF1FFEBFFECFFF3FFFE00090011001400100006FFFBFFF1FFECFFED",
		INIT_70=>X"FFFC00080012001500120009FFFDFFF1FFEBFFEBFFF2FFFD0009001200150011",
		INIT_71=>X"FFFEFFF2FFEAFFE9FFEFFFFB0008001200160013000AFFFDFFF1FFEAFFEAFFF0",
		INIT_72=>X"0006001200180016000DFFFFFFF2FFE9FFE7FFEDFFF90007001200170015000B",
		INIT_73=>X"FFF3FFE7FFE4FFEAFFF600060013001A0018000F0001FFF2FFE8FFE6FFECFFF8",
		INIT_74=>X"0013001C001C00130003FFF3FFE7FFE3FFE8FFF500050013001B001A00110002",
		INIT_75=>X"FFE5FFDFFFE3FFF000020013001E001E00150005FFF3FFE6FFE1FFE6FFF30004",
		INIT_76=>X"00210023001A0009FFF5FFE4FFDDFFE0FFEE00010013001F002100170007FFF4",
		INIT_77=>X"FFD7FFDAFFE8FFFE001400230026001E000BFFF5FFE3FFDAFFDDFFEB00000014",
		INIT_78=>X"002E00260011FFF7FFE1FFD4FFD6FFE4FFFC00140025002A0021000EFFF6FFE2",
		INIT_79=>X"FFCBFFDBFFF60014002B0033002B0015FFF9FFDFFFD0FFD1FFE0FFF900140028",
		INIT_7A=>X"003A0020FFFDFFDBFFC6FFC3FFD4FFF20014002F003A0032001AFFFAFFDDFFCB",
		INIT_7B=>X"FFC0FFE70014003A004B00450028FFFFFFD8FFBEFFBAFFCCFFEE001400330041",
		INIT_7C=>X"00420009FFCFFFA6FF9BFFB1FFDE001400420059005300330003FFD4FFB4FFAD",
		INIT_7D=>X"FFBA00150063008E008A005B0012FFC6FF90FF80FF99FFD10014004F006E0068",
		INIT_7E=>X"0047FF95FF17FEEEFF1CFF8B0015008B00CD00CA00890021FFB7FF6BFF52FF70",
		INIT_7F=>X"0BB80B15094C06B503CB0111FEF6FDBFFD78FDF9FEF8001500FC0175016D00F8",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_10,
		DOPADOP=>dopadop_10,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_11: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"000FFC003FF003FFC00FFF003FFC00FFF003FFC00FFF003FF000FFC003FF000F",
		INITP_01=>X"03FF003FFC00FFF003FFC00FFF003FFC00FFF003FF000FFC003FF000FFC003FF",
		INITP_02=>X"FFC00FFF003FFC00FFF003FFC00FFF003FF000FFC003FF000FFC003FF000FFC0",
		INITP_03=>X"F003FFC00FFF003FFC00FFF003FF000FFC003FF000FFC003FF000FFC003FF003",
		INITP_04=>X"00FFF003FFC00FFF003FF000FFC003FF000FFC003FF000FFC003FF003FFC00FF",
		INITP_05=>X"3FFC00FFF003FF000FFC003FF000FFC003FF000FFC003FF003FFC00FFF003FFC",
		INITP_06=>X"FF003FF000FFC003FF000FFC003FF000FFC003FF003FFC00FFF003FFC00FFF00",
		INITP_07=>X"000FFC003FF000FFC003FF000FFC003FF003FFC00FFF003FFC00FFF003FFC00F",
		INITP_08=>X"F00FF03FC03FC03FC03FC03FC0FF00FF00FF00FF00FF03FC03FC03FC03FC03FC",
		INITP_09=>X"3FC03FC03F00FF00FF00FF00FF00FF03FC03FC03FC03FC03FC0FF00FF00FF00F",
		INITP_0A=>X"00FF00FF00FF00FC03FC03FC03FC03FC03F00FF00FF00FF00FF00FC03FC03FC0",
		INITP_0B=>X"FC03FC03FC03FC03FC03F00FF00FF00FF00FF00FC03FC03FC03FC03FC03F00FF",
		INITP_0C=>X"03FC0FF00FF00FF00FF00FF00FC03FC03FC03FC03FC03F00FF00FF00FF00FF00",
		INITP_0D=>X"F00FF00FF03FC03FC03FC03FC03FC0FF00FF00FF00FF00FF03FC03FC03FC03FC",
		INITP_0E=>X"3FC03FC03FC03FC0FF00FF00FF00FF00FF03FC03FC03FC03FC03FC0FF00FF00F",
		INITP_0F=>X"00FF00FF00FF00FF00FF03FC03FC03FC03FC03FC0FF00FF00FF00FF00FF03FC0",
		INIT_00=>X"000700050001FFFDFFF9FFF8FFF9FFFC000000050007000700050001FFFCFFF9",
		INIT_01=>X"FFF8FFFB000000040007000700050001FFFDFFF9FFF8FFF8FFFC000000040007",
		INIT_02=>X"00060002FFFEFFFAFFF8FFF8FFFBFFFF00040007000700060002FFFDFFF9FFF8",
		INIT_03=>X"FFFAFFFF00030006000800060002FFFEFFFAFFF8FFF8FFFBFFFF000300070007",
		INIT_04=>X"0003FFFFFFFAFFF8FFF8FFFAFFFE00030006000800060003FFFEFFFAFFF8FFF8",
		INIT_05=>X"FFFE00020006000800070003FFFFFFFBFFF8FFF8FFFAFFFE0002000600080006",
		INIT_06=>X"0000FFFBFFF8FFF7FFF9FFFD00020006000800070004FFFFFFFBFFF8FFF8FFFA",
		INIT_07=>X"000100050007000700040000FFFCFFF8FFF7FFF9FFFD00010005000700070004",
		INIT_08=>X"FFFCFFF9FFF7FFF9FFFC000100050007000700050000FFFCFFF8FFF7FFF9FFFC",
		INIT_09=>X"00040007000800050001FFFDFFF9FFF7FFF8FFFC000000050007000700050001",
		INIT_0A=>X"FFF9FFF7FFF8FFFB000000040007000800060002FFFDFFF9FFF7FFF8FFFB0000",
		INIT_0B=>X"0007000800060002FFFEFFF9FFF7FFF8FFFBFFFF00040007000800060002FFFD",
		INIT_0C=>X"FFF7FFF7FFFAFFFF00030007000800060003FFFEFFFAFFF7FFF8FFFAFFFF0004",
		INIT_0D=>X"000800070003FFFFFFFAFFF7FFF7FFFAFFFE00030007000800070003FFFEFFFA",
		INIT_0E=>X"FFF7FFF9FFFD00020006000800070004FFFFFFFAFFF8FFF7FFFAFFFE00030006",
		INIT_0F=>X"000800040000FFFBFFF8FFF7FFF9FFFD00020006000800070004FFFFFFFBFFF8",
		INIT_10=>X"FFF8FFFC000100060008000800050000FFFBFFF8FFF7FFF9FFFD000200060008",
		INIT_11=>X"00050001FFFCFFF8FFF7FFF8FFFC000100050008000800050001FFFCFFF8FFF7",
		INIT_12=>X"FFFB000000050008000800060001FFFCFFF8FFF7FFF8FFFB0000000500080008",
		INIT_13=>X"0002FFFDFFF9FFF7FFF7FFFB000000050008000800060002FFFDFFF8FFF7FFF8",
		INIT_14=>X"FFFF00040008000900070003FFFDFFF9FFF7FFF7FFFAFFFF0004000800090006",
		INIT_15=>X"FFFEFFF9FFF7FFF7FFFAFFFE00040007000900070003FFFEFFF9FFF7FFF7FFFA",
		INIT_16=>X"00030007000900080004FFFFFFFAFFF7FFF6FFF9FFFE00030007000900070003",
		INIT_17=>X"FFFAFFF7FFF6FFF8FFFD00030007000900080004FFFFFFFAFFF7FFF6FFF9FFFE",
		INIT_18=>X"00070009000900050000FFFAFFF7FFF6FFF8FFFD00020007000900080005FFFF",
		INIT_19=>X"FFF7FFF6FFF7FFFC000100060009000900050000FFFBFFF7FFF6FFF8FFFC0002",
		INIT_1A=>X"0009000900060001FFFBFFF7FFF5FFF7FFFB000100060009000900060001FFFB",
		INIT_1B=>X"FFF5FFF6FFFA000000060009000A00070002FFFCFFF7FFF5FFF7FFFB00010006",
		INIT_1C=>X"000A00080003FFFDFFF8FFF5FFF6FFFA000000050009000A00070002FFFCFFF7",
		INIT_1D=>X"FFF5FFF9FFFF00050009000A00080003FFFDFFF8FFF5FFF6FFF9FFFF00050009",
		INIT_1E=>X"00090004FFFEFFF8FFF5FFF5FFF8FFFE00040009000A00080004FFFDFFF8FFF5",
		INIT_1F=>X"FFF8FFFD00040009000B00090005FFFEFFF9FFF5FFF5FFF8FFFE00040009000B",
		INIT_20=>X"0006FFFFFFF9FFF5FFF4FFF7FFFD00030008000B000A0005FFFFFFF9FFF5FFF4",
		INIT_21=>X"FFFB00020008000B000A00060000FFF9FFF5FFF4FFF7FFFC00030008000B000A",
		INIT_22=>X"0001FFFAFFF5FFF3FFF6FFFB00020008000B000B00070000FFFAFFF5FFF4FFF6",
		INIT_23=>X"00010007000B000C00080002FFFBFFF5FFF3FFF5FFFA00010008000B000B0007",
		INIT_24=>X"FFFBFFF5FFF3FFF4FFF900000007000B000C00090002FFFBFFF5FFF3FFF5FFFA",
		INIT_25=>X"0006000C000D000A0003FFFCFFF6FFF2FFF3FFF800000007000C000C00090003",
		INIT_26=>X"FFF6FFF2FFF2FFF7FFFE0006000C000D000A0004FFFCFFF6FFF2FFF3FFF8FFFF",
		INIT_27=>X"000B000E000C0006FFFDFFF6FFF2FFF2FFF6FFFE0006000C000E000B0005FFFD",
		INIT_28=>X"FFF2FFF1FFF5FFFC0005000B000E000C0006FFFEFFF6FFF2FFF1FFF6FFFD0005",
		INIT_29=>X"000F000E0008FFFFFFF7FFF1FFF0FFF4FFFC0004000B000F000D0007FFFFFFF7",
		INIT_2A=>X"FFEFFFF3FFFA0003000B000F000E00090000FFF7FFF1FFF0FFF3FFFB0004000B",
		INIT_2B=>X"0010000A0002FFF8FFF1FFEFFFF2FFF90003000B0010000F000A0001FFF8FFF1",
		INIT_2C=>X"FFF0FFF70001000A00100010000B0002FFF9FFF1FFEEFFF1FFF80002000B0010",
		INIT_2D=>X"000D0004FFFAFFF1FFEDFFEFFFF60000000A00100011000C0003FFF9FFF1FFEE",
		INIT_2E=>X"FFF4FFFF000A00110013000E0005FFFAFFF1FFEDFFEEFFF50000000A00110012",
		INIT_2F=>X"0008FFFCFFF1FFEBFFECFFF3FFFE00090011001400100006FFFBFFF1FFECFFED",
		INIT_30=>X"FFFC00080012001500120009FFFDFFF1FFEBFFEBFFF2FFFD0009001200150011",
		INIT_31=>X"FFFEFFF2FFEAFFE9FFEFFFFB0008001200160013000AFFFDFFF1FFEAFFEAFFF0",
		INIT_32=>X"0006001200180016000DFFFFFFF2FFE9FFE7FFEDFFF90007001200170015000B",
		INIT_33=>X"FFF3FFE7FFE4FFEAFFF600060013001A0018000F0001FFF2FFE8FFE6FFECFFF8",
		INIT_34=>X"0013001C001C00130003FFF3FFE7FFE3FFE8FFF500050013001B001A00110002",
		INIT_35=>X"FFE5FFDFFFE3FFF000020013001E001E00150005FFF3FFE6FFE1FFE6FFF30004",
		INIT_36=>X"00210023001A0009FFF5FFE4FFDDFFE0FFEE00010013001F002100170007FFF4",
		INIT_37=>X"FFD7FFDAFFE8FFFE001400230026001E000BFFF5FFE3FFDAFFDDFFEB00000014",
		INIT_38=>X"002E00260011FFF7FFE1FFD4FFD6FFE4FFFC00140025002A0021000EFFF6FFE2",
		INIT_39=>X"FFCBFFDBFFF60014002B0033002B0015FFF9FFDFFFD0FFD1FFE0FFF900140028",
		INIT_3A=>X"003A0020FFFDFFDBFFC6FFC3FFD4FFF20014002F003A0032001AFFFAFFDDFFCB",
		INIT_3B=>X"FFC0FFE70014003A004B00450028FFFFFFD8FFBEFFBAFFCCFFEE001400330041",
		INIT_3C=>X"00420009FFCFFFA6FF9BFFB1FFDE001400420059005300330003FFD4FFB4FFAD",
		INIT_3D=>X"FFBA00150063008E008A005B0012FFC6FF90FF80FF99FFD10014004F006E0068",
		INIT_3E=>X"0047FF95FF17FEEEFF1CFF8B0015008B00CD00CA00890021FFB7FF6BFF52FF70",
		INIT_3F=>X"0BB80B15094C06B503CB0111FEF6FDBFFD78FDF9FEF8001500FC0175016D00F8",
		INIT_40=>X"000700070002FFFBFFF8FFF9FFFE0004000700060000FFFAFFF8FFFAFFFF0005",
		INIT_41=>X"000600070004FFFEFFF9FFF8FFFC0002000700070003FFFDFFF8FFF8FFFD0003",
		INIT_42=>X"0004000700060000FFFAFFF8FFFAFFFF000500080005FFFFFFF9FFF8FFFA0001",
		INIT_43=>X"0002000700070003FFFDFFF8FFF8FFFD0003000700070002FFFBFFF8FFF9FFFE",
		INIT_44=>X"FFFF000500080005FFFFFFF9FFF7FFFA0001000600070004FFFEFFF9FFF8FFFC",
		INIT_45=>X"FFFD0003000700070002FFFBFFF8FFF9FFFE0004000700060000FFFAFFF7FFFA",
		INIT_46=>X"FFFB0001000600070004FFFEFFF9FFF8FFFC0002000700070003FFFCFFF8FFF8",
		INIT_47=>X"FFF9FFFE0004000800060000FFFAFFF7FFFAFFFF000500080005FFFFFFF9FFF7",
		INIT_48=>X"FFF8FFFC0002000700070003FFFCFFF8FFF8FFFD0003000700070002FFFBFFF8",
		INIT_49=>X"FFF7FFFAFFFF000500080005FFFFFFF9FFF7FFFA0001000600080004FFFEFFF8",
		INIT_4A=>X"FFF8FFF8FFFD0003000700070002FFFBFFF7FFF9FFFE0004000800060000FFFA",
		INIT_4B=>X"FFF9FFF7FFFA0001000600080004FFFEFFF8FFF7FFFC0002000700070003FFFC",
		INIT_4C=>X"FFFBFFF7FFF9FFFE0005000800060000FFFAFFF7FFF9FFFF000600080005FFFF",
		INIT_4D=>X"FFFDFFF8FFF7FFFC0002000700070003FFFCFFF8FFF8FFFD0003000800070002",
		INIT_4E=>X"0000FFFAFFF7FFF90000000600080005FFFFFFF9FFF7FFFA0001000700080004",
		INIT_4F=>X"0003FFFCFFF7FFF8FFFD0004000800070001FFFBFFF7FFF8FFFE000500080006",
		INIT_50=>X"0005FFFFFFF9FFF7FFFA0001000700080004FFFDFFF8FFF7FFFC000200070008",
		INIT_51=>X"00070001FFFBFFF7FFF8FFFE0005000800060000FFFAFFF7FFF9000000060008",
		INIT_52=>X"00080004FFFDFFF8FFF7FFFC0002000800080003FFFCFFF7FFF8FFFD00040008",
		INIT_53=>X"000900060000FFF9FFF6FFF90000000600080005FFFFFFF8FFF7FFFA00010007",
		INIT_54=>X"000800080003FFFCFFF7FFF7FFFD0004000800070001FFFAFFF7FFF8FFFE0005",
		INIT_55=>X"000600090005FFFEFFF8FFF6FFFA0001000700090004FFFDFFF7FFF7FFFB0003",
		INIT_56=>X"0004000900080001FFFAFFF6FFF8FFFE0005000900070000FFF9FFF6FFF90000",
		INIT_57=>X"0001000800090004FFFDFFF7FFF6FFFB0003000800080003FFFBFFF7FFF7FFFD",
		INIT_58=>X"FFFE0006000900070000FFF9FFF6FFF90000000700090006FFFEFFF8FFF6FFFA",
		INIT_59=>X"FFFB0003000900090003FFFBFFF6FFF7FFFD0004000900080001FFFAFFF6FFF8",
		INIT_5A=>X"FFF900000007000A0006FFFEFFF7FFF6FFFA0002000800090004FFFDFFF7FFF6",
		INIT_5B=>X"FFF6FFFD0005000A00080001FFFAFFF5FFF7FFFE0006000A00070000FFF8FFF5",
		INIT_5C=>X"FFF5FFFA00020008000A0005FFFCFFF6FFF6FFFB0003000900090003FFFBFFF6",
		INIT_5D=>X"FFF5FFF7FFFE0006000A00070000FFF8FFF5FFF800000008000A0006FFFEFFF7",
		INIT_5E=>X"FFF6FFF5FFFB0004000A000A0003FFFBFFF5FFF6FFFD0005000A00090002FFF9",
		INIT_5F=>X"FFF8FFF4FFF800000008000B0006FFFEFFF6FFF5FFF900020009000A0005FFFC",
		INIT_60=>X"FFFAFFF4FFF5FFFD0005000B00090002FFF9FFF4FFF7FFFE0007000B00080000",
		INIT_61=>X"FFFEFFF6FFF4FFF90002000A000B0005FFFCFFF5FFF4FFFB0004000A000A0003",
		INIT_62=>X"0002FFF8FFF3FFF6FFFE0007000C00080000FFF7FFF3FFF700000009000B0007",
		INIT_63=>X"0005FFFCFFF4FFF4FFFA0004000B000B0004FFFAFFF4FFF5FFFC0006000C000A",
		INIT_64=>X"00090000FFF6FFF3FFF700000009000C0007FFFEFFF5FFF3FFF90002000A000C",
		INIT_65=>X"000C0004FFF9FFF3FFF4FFFC0007000C000A0002FFF8FFF2FFF5FFFE0008000D",
		INIT_66=>X"000D0008FFFDFFF4FFF2FFF80003000B000D0006FFFBFFF3FFF3FFFA0005000C",
		INIT_67=>X"000E000B0002FFF7FFF1FFF5FFFE0009000E000AFFFFFFF5FFF1FFF60001000A",
		INIT_68=>X"000D000E0006FFFBFFF2FFF2FFFA0005000D000D0004FFF9FFF2FFF3FFFC0007",
		INIT_69=>X"000A000F000BFFFFFFF4FFF0FFF50001000B000F0009FFFDFFF3FFF1FFF80003",
		INIT_6A=>X"0006000F000E0004FFF8FFF0FFF2FFFC0008000F000C0002FFF6FFF0FFF4FFFE",
		INIT_6B=>X"0001000D00100009FFFDFFF2FFEFFFF70004000E000F0007FFFAFFF1FFF0FFF9",
		INIT_6C=>X"FFFC00090011000E0002FFF5FFEEFFF2FFFE000B0011000CFFFFFFF3FFEEFFF4",
		INIT_6D=>X"FFF60004001000110008FFF9FFEFFFEFFFF90007001100100005FFF7FFEEFFF0",
		INIT_6E=>X"FFF1FFFE000D0013000DFFFFFFF1FFECFFF30002000F0012000BFFFCFFF0FFED",
		INIT_6F=>X"FFECFFF80008001300120005FFF5FFECFFEEFFFB000B001300100002FFF3FFEC",
		INIT_70=>X"FFE9FFF1000200110015000CFFFBFFEDFFEBFFF50005001200140009FFF8FFEC",
		INIT_71=>X"FFE8FFEBFFFB000D001700120002FFF1FFE9FFEEFFFE000F0016000FFFFFFFEF",
		INIT_72=>X"FFEAFFE7FFF3000600160017000AFFF7FFE9FFE9FFF7000A001600150006FFF4",
		INIT_73=>X"FFEEFFE4FFEBFFFE0012001A0012FFFEFFECFFE5FFEF000300140019000EFFFA",
		INIT_74=>X"FFF5FFE4FFE4FFF5000C001B00190007FFF1FFE4FFE8FFFA0010001B00160003",
		INIT_75=>X"FFFEFFE7FFDFFFEB00040019001F0011FFF9FFE5FFE1FFF00008001B001C000C",
		INIT_76=>X"0009FFEDFFDCFFE1FFF900140022001B0003FFE9FFDDFFE6FFFE001700210016",
		INIT_77=>X"0016FFF7FFDDFFD9FFEC000B002200240010FFF1FFDCFFDDFFF3001000230020",
		INIT_78=>X"00240004FFE2FFD2FFDEFFFE001F002C001DFFFDFFDFFFD5FFE5000500210028",
		INIT_79=>X"00330016FFECFFCEFFD0FFEE00160030002C000CFFE6FFD0FFD7FFF7001B002E",
		INIT_7A=>X"0041002BFFFBFFCFFFC2FFDA00080030003A0020FFF3FFCEFFC9FFE400100031",
		INIT_7B=>X"004E00460013FFD7FFB4FFC1FFF3002B004700380006FFD2FFBBFFCEFFFE002F",
		INIT_7C=>X"005800680038FFE8FFA9FFA1FFD2001D005300560024FFDEFFAEFFB2FFE40025",
		INIT_7D=>X"0061009C0077000DFFA0FF73FF9CFFFE005D007F0053FFF7FFA4FF8CFFBB0010",
		INIT_7E=>X"00660114010F006CFF9AFF18FF29FFB7006400C800AE002FFF9DFF4FFF70FFE3",
		INIT_7F=>X"10680EB00A2D0481FF98FCD8FCA1FE3F006701DC01FF00FEFF98FEA5FE99FF5D",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_11,
		DOPADOP=>dopadop_11,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_12: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"F00FF03FC03FC03FC03FC03FC0FF00FF00FF00FF00FF03FC03FC03FC03FC03FC",
		INITP_01=>X"3FC03FC03F00FF00FF00FF00FF00FF03FC03FC03FC03FC03FC0FF00FF00FF00F",
		INITP_02=>X"00FF00FF00FF00FC03FC03FC03FC03FC03F00FF00FF00FF00FF00FC03FC03FC0",
		INITP_03=>X"FC03FC03FC03FC03FC03F00FF00FF00FF00FF00FC03FC03FC03FC03FC03F00FF",
		INITP_04=>X"03FC0FF00FF00FF00FF00FF00FC03FC03FC03FC03FC03F00FF00FF00FF00FF00",
		INITP_05=>X"F00FF00FF03FC03FC03FC03FC03FC0FF00FF00FF00FF00FF03FC03FC03FC03FC",
		INITP_06=>X"3FC03FC03FC03FC0FF00FF00FF00FF00FF03FC03FC03FC03FC03FC0FF00FF00F",
		INITP_07=>X"00FF00FF00FF00FF00FF03FC03FC03FC03FC03FC0FF00FF00FF00FF00FF03FC0",
		INITP_08=>X"F03C0FC0F03F03F0FC0FC0F03F03C0FC0FC3F03F03C0FC0F03F03F0FC0FC0F03",
		INITP_09=>X"F0FC0FC3F03F03C0FC0FC3F03F0FC0FC0F03F03F0FC0FC3F03F03C0FC0FC3F03",
		INITP_0A=>X"C0FC0FC3F03F0FC0FC0F03F03F0FC0FC3F03F03C0FC0FC3F03F0FC0FC0F03F03",
		INITP_0B=>X"C0FC0F03F03C0FC0FC3F03F03C0FC0F03F03F0FC0FC0F03F03F0FC0FC3F03F03",
		INITP_0C=>X"C0FC3F03F03C0FC0F03F03F0FC0FC0F03F03C0FC0FC3F03F03C0FC0F03F03F0F",
		INITP_0D=>X"C0F03F03F0FC0FC3F03F03C0FC0FC3F03F03C0FC0F03F03F0FC0FC0F03F03C0F",
		INITP_0E=>X"C3F03F03C0FC0FC3F03F0FC0FC0F03F03F0FC0FC3F03F03C0FC0FC3F03F0FC0F",
		INITP_0F=>X"03F03F0FC0FC0F03F03F0FC0FC3F03F03C0FC0FC3F03F0FC0FC0F03F03F0FC0F",
		INIT_00=>X"000700070002FFFBFFF8FFF9FFFE0004000700060000FFFAFFF8FFFAFFFF0005",
		INIT_01=>X"000600070004FFFEFFF9FFF8FFFC0002000700070003FFFDFFF8FFF8FFFD0003",
		INIT_02=>X"0004000700060000FFFAFFF8FFFAFFFF000500080005FFFFFFF9FFF8FFFA0001",
		INIT_03=>X"0002000700070003FFFDFFF8FFF8FFFD0003000700070002FFFBFFF8FFF9FFFE",
		INIT_04=>X"FFFF000500080005FFFFFFF9FFF7FFFA0001000600070004FFFEFFF9FFF8FFFC",
		INIT_05=>X"FFFD0003000700070002FFFBFFF8FFF9FFFE0004000700060000FFFAFFF7FFFA",
		INIT_06=>X"FFFB0001000600070004FFFEFFF9FFF8FFFC0002000700070003FFFCFFF8FFF8",
		INIT_07=>X"FFF9FFFE0004000800060000FFFAFFF7FFFAFFFF000500080005FFFFFFF9FFF7",
		INIT_08=>X"FFF8FFFC0002000700070003FFFCFFF8FFF8FFFD0003000700070002FFFBFFF8",
		INIT_09=>X"FFF7FFFAFFFF000500080005FFFFFFF9FFF7FFFA0001000600080004FFFEFFF8",
		INIT_0A=>X"FFF8FFF8FFFD0003000700070002FFFBFFF7FFF9FFFE0004000800060000FFFA",
		INIT_0B=>X"FFF9FFF7FFFA0001000600080004FFFEFFF8FFF7FFFC0002000700070003FFFC",
		INIT_0C=>X"FFFBFFF7FFF9FFFE0005000800060000FFFAFFF7FFF9FFFF000600080005FFFF",
		INIT_0D=>X"FFFDFFF8FFF7FFFC0002000700070003FFFCFFF8FFF8FFFD0003000800070002",
		INIT_0E=>X"0000FFFAFFF7FFF90000000600080005FFFFFFF9FFF7FFFA0001000700080004",
		INIT_0F=>X"0003FFFCFFF7FFF8FFFD0004000800070001FFFBFFF7FFF8FFFE000500080006",
		INIT_10=>X"0005FFFFFFF9FFF7FFFA0001000700080004FFFDFFF8FFF7FFFC000200070008",
		INIT_11=>X"00070001FFFBFFF7FFF8FFFE0005000800060000FFFAFFF7FFF9000000060008",
		INIT_12=>X"00080004FFFDFFF8FFF7FFFC0002000800080003FFFCFFF7FFF8FFFD00040008",
		INIT_13=>X"000900060000FFF9FFF6FFF90000000600080005FFFFFFF8FFF7FFFA00010007",
		INIT_14=>X"000800080003FFFCFFF7FFF7FFFD0004000800070001FFFAFFF7FFF8FFFE0005",
		INIT_15=>X"000600090005FFFEFFF8FFF6FFFA0001000700090004FFFDFFF7FFF7FFFB0003",
		INIT_16=>X"0004000900080001FFFAFFF6FFF8FFFE0005000900070000FFF9FFF6FFF90000",
		INIT_17=>X"0001000800090004FFFDFFF7FFF6FFFB0003000800080003FFFBFFF7FFF7FFFD",
		INIT_18=>X"FFFE0006000900070000FFF9FFF6FFF90000000700090006FFFEFFF8FFF6FFFA",
		INIT_19=>X"FFFB0003000900090003FFFBFFF6FFF7FFFD0004000900080001FFFAFFF6FFF8",
		INIT_1A=>X"FFF900000007000A0006FFFEFFF7FFF6FFFA0002000800090004FFFDFFF7FFF6",
		INIT_1B=>X"FFF6FFFD0005000A00080001FFFAFFF5FFF7FFFE0006000A00070000FFF8FFF5",
		INIT_1C=>X"FFF5FFFA00020008000A0005FFFCFFF6FFF6FFFB0003000900090003FFFBFFF6",
		INIT_1D=>X"FFF5FFF7FFFE0006000A00070000FFF8FFF5FFF800000008000A0006FFFEFFF7",
		INIT_1E=>X"FFF6FFF5FFFB0004000A000A0003FFFBFFF5FFF6FFFD0005000A00090002FFF9",
		INIT_1F=>X"FFF8FFF4FFF800000008000B0006FFFEFFF6FFF5FFF900020009000A0005FFFC",
		INIT_20=>X"FFFAFFF4FFF5FFFD0005000B00090002FFF9FFF4FFF7FFFE0007000B00080000",
		INIT_21=>X"FFFEFFF6FFF4FFF90002000A000B0005FFFCFFF5FFF4FFFB0004000A000A0003",
		INIT_22=>X"0002FFF8FFF3FFF6FFFE0007000C00080000FFF7FFF3FFF700000009000B0007",
		INIT_23=>X"0005FFFCFFF4FFF4FFFA0004000B000B0004FFFAFFF4FFF5FFFC0006000C000A",
		INIT_24=>X"00090000FFF6FFF3FFF700000009000C0007FFFEFFF5FFF3FFF90002000A000C",
		INIT_25=>X"000C0004FFF9FFF3FFF4FFFC0007000C000A0002FFF8FFF2FFF5FFFE0008000D",
		INIT_26=>X"000D0008FFFDFFF4FFF2FFF80003000B000D0006FFFBFFF3FFF3FFFA0005000C",
		INIT_27=>X"000E000B0002FFF7FFF1FFF5FFFE0009000E000AFFFFFFF5FFF1FFF60001000A",
		INIT_28=>X"000D000E0006FFFBFFF2FFF2FFFA0005000D000D0004FFF9FFF2FFF3FFFC0007",
		INIT_29=>X"000A000F000BFFFFFFF4FFF0FFF50001000B000F0009FFFDFFF3FFF1FFF80003",
		INIT_2A=>X"0006000F000E0004FFF8FFF0FFF2FFFC0008000F000C0002FFF6FFF0FFF4FFFE",
		INIT_2B=>X"0001000D00100009FFFDFFF2FFEFFFF70004000E000F0007FFFAFFF1FFF0FFF9",
		INIT_2C=>X"FFFC00090011000E0002FFF5FFEEFFF2FFFE000B0011000CFFFFFFF3FFEEFFF4",
		INIT_2D=>X"FFF60004001000110008FFF9FFEFFFEFFFF90007001100100005FFF7FFEEFFF0",
		INIT_2E=>X"FFF1FFFE000D0013000DFFFFFFF1FFECFFF30002000F0012000BFFFCFFF0FFED",
		INIT_2F=>X"FFECFFF80008001300120005FFF5FFECFFEEFFFB000B001300100002FFF3FFEC",
		INIT_30=>X"FFE9FFF1000200110015000CFFFBFFEDFFEBFFF50005001200140009FFF8FFEC",
		INIT_31=>X"FFE8FFEBFFFB000D001700120002FFF1FFE9FFEEFFFE000F0016000FFFFFFFEF",
		INIT_32=>X"FFEAFFE7FFF3000600160017000AFFF7FFE9FFE9FFF7000A001600150006FFF4",
		INIT_33=>X"FFEEFFE4FFEBFFFE0012001A0012FFFEFFECFFE5FFEF000300140019000EFFFA",
		INIT_34=>X"FFF5FFE4FFE4FFF5000C001B00190007FFF1FFE4FFE8FFFA0010001B00160003",
		INIT_35=>X"FFFEFFE7FFDFFFEB00040019001F0011FFF9FFE5FFE1FFF00008001B001C000C",
		INIT_36=>X"0009FFEDFFDCFFE1FFF900140022001B0003FFE9FFDDFFE6FFFE001700210016",
		INIT_37=>X"0016FFF7FFDDFFD9FFEC000B002200240010FFF1FFDCFFDDFFF3001000230020",
		INIT_38=>X"00240004FFE2FFD2FFDEFFFE001F002C001DFFFDFFDFFFD5FFE5000500210028",
		INIT_39=>X"00330016FFECFFCEFFD0FFEE00160030002C000CFFE6FFD0FFD7FFF7001B002E",
		INIT_3A=>X"0041002BFFFBFFCFFFC2FFDA00080030003A0020FFF3FFCEFFC9FFE400100031",
		INIT_3B=>X"004E00460013FFD7FFB4FFC1FFF3002B004700380006FFD2FFBBFFCEFFFE002F",
		INIT_3C=>X"005800680038FFE8FFA9FFA1FFD2001D005300560024FFDEFFAEFFB2FFE40025",
		INIT_3D=>X"0061009C0077000DFFA0FF73FF9CFFFE005D007F0053FFF7FFA4FF8CFFBB0010",
		INIT_3E=>X"00660114010F006CFF9AFF18FF29FFB7006400C800AE002FFF9DFF4FFF70FFE3",
		INIT_3F=>X"10680EB00A2D0481FF98FCD8FCA1FE3F006701DC01FF00FEFF98FEA5FE99FF5D",
		INIT_40=>X"FFFA000200070003FFFBFFF8FFFD000600070000FFF8FFF9000100070005FFFC",
		INIT_41=>X"000000070005FFFDFFF8FFFB000400070002FFFAFFF8FFFF00060006FFFEFFF8",
		INIT_42=>X"000600070000FFF8FFF9000100070004FFFCFFF7FFFC000500070001FFF9FFF8",
		INIT_43=>X"00080002FFFAFFF8FFFF00060006FFFEFFF8FFFA000200080003FFFBFFF8FFFD",
		INIT_44=>X"0004FFFCFFF7FFFC000500070001FFF9FFF8000000070005FFFDFFF8FFFB0004",
		INIT_45=>X"FFFEFFF8FFFA000300080003FFFBFFF8FFFD000600070000FFF8FFF900010007",
		INIT_46=>X"FFF9FFF8000000070005FFFDFFF7FFFB000400080002FFFAFFF8FFFF00060006",
		INIT_47=>X"FFF8FFFE000600070000FFF8FFF9000100070004FFFCFFF7FFFC000500070001",
		INIT_48=>X"FFFB000400080002FFFAFFF8FFFF00070006FFFEFFF8FFFA000300080003FFFB",
		INIT_49=>X"000200080004FFFCFFF7FFFC000500070001FFF9FFF8000000070005FFFDFFF7",
		INIT_4A=>X"00070006FFFEFFF8FFFA000300080003FFFAFFF7FFFE00060007FFFFFFF8FFF9",
		INIT_4B=>X"00080001FFF9FFF8000000070005FFFDFFF7FFFB000400080002FFF9FFF8FFFF",
		INIT_4C=>X"0003FFFAFFF7FFFE00060007FFFFFFF8FFF9000200080004FFFCFFF7FFFC0005",
		INIT_4D=>X"FFFDFFF7FFFB000400080002FFF9FFF8FFFF00070006FFFEFFF7FFFA00030008",
		INIT_4E=>X"FFF8FFF9000200080004FFFBFFF7FFFC000500080001FFF8FFF8000000080006",
		INIT_4F=>X"FFF8FFFF00070006FFFEFFF7FFFA000300080003FFFAFFF7FFFE00060007FFFF",
		INIT_50=>X"FFFC000600080001FFF8FFF8000000080006FFFCFFF7FFFB000400080002FFF9",
		INIT_51=>X"000300080003FFFAFFF7FFFE00070007FFFFFFF7FFF9000200080005FFFBFFF7",
		INIT_52=>X"00080006FFFCFFF7FFFB000500080002FFF9FFF7FFFF00070007FFFEFFF7FFFA",
		INIT_53=>X"0008FFFFFFF7FFF9000200080005FFFBFFF7FFFC000600080001FFF8FFF80001",
		INIT_54=>X"0002FFF9FFF7FFFF00080007FFFEFFF7FFFA000300090003FFFAFFF7FFFE0007",
		INIT_55=>X"FFFBFFF6FFFC000600080000FFF8FFF8000100080006FFFCFFF6FFFB00050009",
		INIT_56=>X"FFF6FFFA000400090003FFF9FFF6FFFE00070008FFFFFFF7FFF9000200090005",
		INIT_57=>X"FFF8000100090006FFFCFFF6FFFB000500090002FFF8FFF7FFFF00080007FFFD",
		INIT_58=>X"FFFE00070008FFFFFFF6FFF8000200090005FFFAFFF6FFFC000600090000FFF7",
		INIT_59=>X"000500090002FFF8FFF7FFFF00080007FFFDFFF6FFFA000400090003FFF9FFF6",
		INIT_5A=>X"000A0005FFFAFFF5FFFC000700090000FFF7FFF7000100090006FFFCFFF6FFFB",
		INIT_5B=>X"0008FFFDFFF5FFF90004000A0004FFF9FFF6FFFE00080008FFFFFFF6FFF80003",
		INIT_5C=>X"0000FFF6FFF70001000A0006FFFBFFF5FFFB0006000A0002FFF7FFF600000009",
		INIT_5D=>X"FFF8FFF5FFFE00080009FFFFFFF5FFF80003000A0005FFFAFFF5FFFC00070009",
		INIT_5E=>X"FFF4FFFB0006000A0002FFF7FFF6000000090008FFFDFFF5FFF90005000A0004",
		INIT_5F=>X"FFF80003000B0005FFF9FFF4FFFC0008000A0000FFF6FFF60001000A0007FFFB",
		INIT_60=>X"0000000A0008FFFCFFF4FFF90005000B0004FFF8FFF5FFFE00090009FFFEFFF5",
		INIT_61=>X"0008000A0000FFF5FFF60002000B0007FFFBFFF4FFFA0007000B0002FFF6FFF5",
		INIT_62=>X"000C0004FFF7FFF4FFFE000A000AFFFEFFF4FFF70004000B0006FFF9FFF4FFFC",
		INIT_63=>X"0008FFFAFFF3FFFA0007000C0002FFF6FFF40000000B0009FFFCFFF3FFF80006",
		INIT_64=>X"FFFEFFF3FFF70004000C0006FFF8FFF3FFFC0009000B0000FFF4FFF50002000C",
		INIT_65=>X"FFF5FFF40000000C0009FFFCFFF2FFF80006000D0004FFF6FFF3FFFE000B000A",
		INIT_66=>X"FFF2FFFC000A000C0000FFF3FFF50002000D0008FFFAFFF2FFFA0008000D0002",
		INIT_67=>X"FFF80007000E0004FFF5FFF2FFFE000C000BFFFEFFF2FFF60005000D0006FFF7",
		INIT_68=>X"0003000E0009FFF9FFF1FFF90009000E0002FFF4FFF30000000D000AFFFBFFF1",
		INIT_69=>X"000D000CFFFDFFF1FFF50005000F0007FFF7FFF1FFFC000B000D0000FFF2FFF4",
		INIT_6A=>X"000F0002FFF2FFF10001000E000BFFFBFFF0FFF70008000F0005FFF4FFF1FFFE",
		INIT_6B=>X"0008FFF5FFEFFFFB000C000F0000FFF1FFF300030010000AFFF8FFEFFFF9000A",
		INIT_6C=>X"FFFAFFEEFFF6000900110005FFF3FFEFFFFE000E000EFFFDFFEFFFF400060011",
		INIT_6D=>X"FFEFFFF100040012000BFFF7FFEDFFF8000C00110002FFF1FFF000010010000C",
		INIT_6E=>X"FFEDFFFE00110010FFFCFFEDFFF3000700130008FFF4FFEDFFFB000E0011FFFF",
		INIT_6F=>X"FFF8000D00130003FFEEFFEE00010013000EFFF9FFEBFFF5000A00130006FFF1",
		INIT_70=>X"000900160009FFF2FFEAFFFB00100013FFFFFFECFFEF00050014000CFFF6FFEB",
		INIT_71=>X"00160010FFF8FFE8FFF3000C00160006FFEFFFEAFFFE00130012FFFCFFEAFFF1",
		INIT_72=>X"0016FFFFFFE8FFEC00060018000EFFF4FFE7FFF6001000170003FFEBFFEB0002",
		INIT_73=>X"0008FFEBFFE6FFFE00170015FFFBFFE6FFEE000A001A000BFFEFFFE6FFFA0014",
		INIT_74=>X"FFF1FFE2FFF50014001B0003FFE7FFE70003001B0013FFF6FFE3FFF1000F001B",
		INIT_75=>X"FFE0FFEB000D0020000DFFEBFFE1FFF90018001BFFFEFFE3FFE80008001D0011",
		INIT_76=>X"FFE1000400220018FFF3FFDCFFEE001300220009FFE6FFE0FFFE001D001AFFF9",
		INIT_77=>X"FFF800200023FFFEFFDBFFE2000B00260015FFECFFDAFFF2001A00230004FFE0",
		INIT_78=>X"001A002D000CFFDDFFD6FFFE00270023FFF6FFD5FFE50012002A0011FFE5FFD7",
		INIT_79=>X"0035001EFFE4FFCBFFEE002400300005FFD5FFD60006002E0021FFEEFFD0FFE8",
		INIT_7A=>X"0033FFF1FFC1FFD9001B003D0019FFD9FFC6FFF5002F0032FFFCFFCBFFD60010",
		INIT_7B=>X"0008FFBBFFBE000B00490033FFE4FFB6FFDD002900450012FFCBFFC2FFFE003B",
		INIT_7C=>X"FFB8FF99FFED00530057FFF9FFA6FFBA001C005A0031FFD1FFA9FFE3003B004E",
		INIT_7D=>X"FF5DFFB5005B00920024FF93FF83FFFE00750063FFE3FF89FFB700340071002C",
		INIT_7E=>X"FF13005F011F0093FF75FF09FFB300A200CB0012FF52FF60001C00AC0074FFBF",
		INIT_7F=>X"16F8126707E4FE61FB02FD8C019202E80100FE80FE0AFFB20164015CFFE3FEBB",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_12,
		DOPADOP=>dopadop_12,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_13: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"F03C0FC0F03F03F0FC0FC0F03F03C0FC0FC3F03F03C0FC0F03F03F0FC0FC0F03",
		INITP_01=>X"F0FC0FC3F03F03C0FC0FC3F03F0FC0FC0F03F03F0FC0FC3F03F03C0FC0FC3F03",
		INITP_02=>X"C0FC0FC3F03F0FC0FC0F03F03F0FC0FC3F03F03C0FC0FC3F03F0FC0FC0F03F03",
		INITP_03=>X"C0FC0F03F03C0FC0FC3F03F03C0FC0F03F03F0FC0FC0F03F03F0FC0FC3F03F03",
		INITP_04=>X"C0FC3F03F03C0FC0F03F03F0FC0FC0F03F03C0FC0FC3F03F03C0FC0F03F03F0F",
		INITP_05=>X"C0F03F03F0FC0FC3F03F03C0FC0FC3F03F03C0FC0F03F03F0FC0FC0F03F03C0F",
		INITP_06=>X"C3F03F03C0FC0FC3F03F0FC0FC0F03F03F0FC0FC3F03F03C0FC0FC3F03F0FC0F",
		INITP_07=>X"03F03F0FC0FC0F03F03F0FC0FC3F03F03C0FC0FC3F03F0FC0FC0F03F03F0FC0F",
		INITP_08=>X"F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0",
		INITP_09=>X"3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C30F0F0F0F0",
		INITP_0A=>X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F3C3C3C3C3C3C3C3C3C",
		INITP_0B=>X"C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3CF0F0F0F0F0F0F0F0F0F0F0F0F0F",
		INITP_0C=>X"F0F0F0F0F0F0F0F0F0F0F0F0F0F3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3",
		INITP_0D=>X"3C3C3C3C3C3C3C3C3C30F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0",
		INITP_0E=>X"0F0F0F0F0C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C",
		INITP_0F=>X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F",
		INIT_00=>X"FFFA000200070003FFFBFFF8FFFD000600070000FFF8FFF9000100070005FFFC",
		INIT_01=>X"000000070005FFFDFFF8FFFB000400070002FFFAFFF8FFFF00060006FFFEFFF8",
		INIT_02=>X"000600070000FFF8FFF9000100070004FFFCFFF7FFFC000500070001FFF9FFF8",
		INIT_03=>X"00080002FFFAFFF8FFFF00060006FFFEFFF8FFFA000200080003FFFBFFF8FFFD",
		INIT_04=>X"0004FFFCFFF7FFFC000500070001FFF9FFF8000000070005FFFDFFF8FFFB0004",
		INIT_05=>X"FFFEFFF8FFFA000300080003FFFBFFF8FFFD000600070000FFF8FFF900010007",
		INIT_06=>X"FFF9FFF8000000070005FFFDFFF7FFFB000400080002FFFAFFF8FFFF00060006",
		INIT_07=>X"FFF8FFFE000600070000FFF8FFF9000100070004FFFCFFF7FFFC000500070001",
		INIT_08=>X"FFFB000400080002FFFAFFF8FFFF00070006FFFEFFF8FFFA000300080003FFFB",
		INIT_09=>X"000200080004FFFCFFF7FFFC000500070001FFF9FFF8000000070005FFFDFFF7",
		INIT_0A=>X"00070006FFFEFFF8FFFA000300080003FFFAFFF7FFFE00060007FFFFFFF8FFF9",
		INIT_0B=>X"00080001FFF9FFF8000000070005FFFDFFF7FFFB000400080002FFF9FFF8FFFF",
		INIT_0C=>X"0003FFFAFFF7FFFE00060007FFFFFFF8FFF9000200080004FFFCFFF7FFFC0005",
		INIT_0D=>X"FFFDFFF7FFFB000400080002FFF9FFF8FFFF00070006FFFEFFF7FFFA00030008",
		INIT_0E=>X"FFF8FFF9000200080004FFFBFFF7FFFC000500080001FFF8FFF8000000080006",
		INIT_0F=>X"FFF8FFFF00070006FFFEFFF7FFFA000300080003FFFAFFF7FFFE00060007FFFF",
		INIT_10=>X"FFFC000600080001FFF8FFF8000000080006FFFCFFF7FFFB000400080002FFF9",
		INIT_11=>X"000300080003FFFAFFF7FFFE00070007FFFFFFF7FFF9000200080005FFFBFFF7",
		INIT_12=>X"00080006FFFCFFF7FFFB000500080002FFF9FFF7FFFF00070007FFFEFFF7FFFA",
		INIT_13=>X"0008FFFFFFF7FFF9000200080005FFFBFFF7FFFC000600080001FFF8FFF80001",
		INIT_14=>X"0002FFF9FFF7FFFF00080007FFFEFFF7FFFA000300090003FFFAFFF7FFFE0007",
		INIT_15=>X"FFFBFFF6FFFC000600080000FFF8FFF8000100080006FFFCFFF6FFFB00050009",
		INIT_16=>X"FFF6FFFA000400090003FFF9FFF6FFFE00070008FFFFFFF7FFF9000200090005",
		INIT_17=>X"FFF8000100090006FFFCFFF6FFFB000500090002FFF8FFF7FFFF00080007FFFD",
		INIT_18=>X"FFFE00070008FFFFFFF6FFF8000200090005FFFAFFF6FFFC000600090000FFF7",
		INIT_19=>X"000500090002FFF8FFF7FFFF00080007FFFDFFF6FFFA000400090003FFF9FFF6",
		INIT_1A=>X"000A0005FFFAFFF5FFFC000700090000FFF7FFF7000100090006FFFCFFF6FFFB",
		INIT_1B=>X"0008FFFDFFF5FFF90004000A0004FFF9FFF6FFFE00080008FFFFFFF6FFF80003",
		INIT_1C=>X"0000FFF6FFF70001000A0006FFFBFFF5FFFB0006000A0002FFF7FFF600000009",
		INIT_1D=>X"FFF8FFF5FFFE00080009FFFFFFF5FFF80003000A0005FFFAFFF5FFFC00070009",
		INIT_1E=>X"FFF4FFFB0006000A0002FFF7FFF6000000090008FFFDFFF5FFF90005000A0004",
		INIT_1F=>X"FFF80003000B0005FFF9FFF4FFFC0008000A0000FFF6FFF60001000A0007FFFB",
		INIT_20=>X"0000000A0008FFFCFFF4FFF90005000B0004FFF8FFF5FFFE00090009FFFEFFF5",
		INIT_21=>X"0008000A0000FFF5FFF60002000B0007FFFBFFF4FFFA0007000B0002FFF6FFF5",
		INIT_22=>X"000C0004FFF7FFF4FFFE000A000AFFFEFFF4FFF70004000B0006FFF9FFF4FFFC",
		INIT_23=>X"0008FFFAFFF3FFFA0007000C0002FFF6FFF40000000B0009FFFCFFF3FFF80006",
		INIT_24=>X"FFFEFFF3FFF70004000C0006FFF8FFF3FFFC0009000B0000FFF4FFF50002000C",
		INIT_25=>X"FFF5FFF40000000C0009FFFCFFF2FFF80006000D0004FFF6FFF3FFFE000B000A",
		INIT_26=>X"FFF2FFFC000A000C0000FFF3FFF50002000D0008FFFAFFF2FFFA0008000D0002",
		INIT_27=>X"FFF80007000E0004FFF5FFF2FFFE000C000BFFFEFFF2FFF60005000D0006FFF7",
		INIT_28=>X"0003000E0009FFF9FFF1FFF90009000E0002FFF4FFF30000000D000AFFFBFFF1",
		INIT_29=>X"000D000CFFFDFFF1FFF50005000F0007FFF7FFF1FFFC000B000D0000FFF2FFF4",
		INIT_2A=>X"000F0002FFF2FFF10001000E000BFFFBFFF0FFF70008000F0005FFF4FFF1FFFE",
		INIT_2B=>X"0008FFF5FFEFFFFB000C000F0000FFF1FFF300030010000AFFF8FFEFFFF9000A",
		INIT_2C=>X"FFFAFFEEFFF6000900110005FFF3FFEFFFFE000E000EFFFDFFEFFFF400060011",
		INIT_2D=>X"FFEFFFF100040012000BFFF7FFEDFFF8000C00110002FFF1FFF000010010000C",
		INIT_2E=>X"FFEDFFFE00110010FFFCFFEDFFF3000700130008FFF4FFEDFFFB000E0011FFFF",
		INIT_2F=>X"FFF8000D00130003FFEEFFEE00010013000EFFF9FFEBFFF5000A00130006FFF1",
		INIT_30=>X"000900160009FFF2FFEAFFFB00100013FFFFFFECFFEF00050014000CFFF6FFEB",
		INIT_31=>X"00160010FFF8FFE8FFF3000C00160006FFEFFFEAFFFE00130012FFFCFFEAFFF1",
		INIT_32=>X"0016FFFFFFE8FFEC00060018000EFFF4FFE7FFF6001000170003FFEBFFEB0002",
		INIT_33=>X"0008FFEBFFE6FFFE00170015FFFBFFE6FFEE000A001A000BFFEFFFE6FFFA0014",
		INIT_34=>X"FFF1FFE2FFF50014001B0003FFE7FFE70003001B0013FFF6FFE3FFF1000F001B",
		INIT_35=>X"FFE0FFEB000D0020000DFFEBFFE1FFF90018001BFFFEFFE3FFE80008001D0011",
		INIT_36=>X"FFE1000400220018FFF3FFDCFFEE001300220009FFE6FFE0FFFE001D001AFFF9",
		INIT_37=>X"FFF800200023FFFEFFDBFFE2000B00260015FFECFFDAFFF2001A00230004FFE0",
		INIT_38=>X"001A002D000CFFDDFFD6FFFE00270023FFF6FFD5FFE50012002A0011FFE5FFD7",
		INIT_39=>X"0035001EFFE4FFCBFFEE002400300005FFD5FFD60006002E0021FFEEFFD0FFE8",
		INIT_3A=>X"0033FFF1FFC1FFD9001B003D0019FFD9FFC6FFF5002F0032FFFCFFCBFFD60010",
		INIT_3B=>X"0008FFBBFFBE000B00490033FFE4FFB6FFDD002900450012FFCBFFC2FFFE003B",
		INIT_3C=>X"FFB8FF99FFED00530057FFF9FFA6FFBA001C005A0031FFD1FFA9FFE3003B004E",
		INIT_3D=>X"FF5DFFB5005B00920024FF93FF83FFFE00750063FFE3FF89FFB700340071002C",
		INIT_3E=>X"FF13005F011F0093FF75FF09FFB300A200CB0012FF52FF60001C00AC0074FFBF",
		INIT_3F=>X"16F8126707E4FE61FB02FD8C019202E80100FE80FE0AFFB20164015CFFE3FEBB",
		INIT_40=>X"FFF8FFFE00070001FFF8FFFF00070000FFF8FFFF00070000FFF8FFFF00070000",
		INIT_41=>X"FFF8FFFD00070002FFF8FFFD00070002FFF8FFFE00070001FFF8FFFE00070001",
		INIT_42=>X"FFF9FFFC00070003FFF8FFFC00070003FFF8FFFC00070003FFF8FFFD00070002",
		INIT_43=>X"FFF9FFFA00060004FFF9FFFB00060004FFF9FFFB00060004FFF9FFFB00060004",
		INIT_44=>X"FFFAFFF900050005FFFAFFFA00050005FFFAFFFA00050005FFFAFFFA00060005",
		INIT_45=>X"FFFBFFF900040006FFFBFFF900040006FFFBFFF900040006FFFAFFF900050006",
		INIT_46=>X"FFFDFFF800030007FFFCFFF800030007FFFCFFF800030007FFFCFFF800040006",
		INIT_47=>X"FFFEFFF800010007FFFEFFF800020007FFFDFFF800020007FFFDFFF800020007",
		INIT_48=>X"FFFFFFF700000008FFFFFFF700000008FFFFFFF700010008FFFEFFF700010008",
		INIT_49=>X"0001FFF7FFFE00080000FFF7FFFF00080000FFF7FFFF00080000FFF700000008",
		INIT_4A=>X"0002FFF8FFFD00070002FFF8FFFD00080001FFF7FFFE00080001FFF7FFFE0008",
		INIT_4B=>X"0003FFF8FFFC00070003FFF8FFFC00070003FFF8FFFC00070002FFF8FFFD0007",
		INIT_4C=>X"0005FFF9FFFA00060004FFF9FFFB00060004FFF8FFFB00070004FFF8FFFB0007",
		INIT_4D=>X"0006FFFAFFF900050006FFF9FFFA00060005FFF9FFFA00060005FFF9FFFA0006",
		INIT_4E=>X"0007FFFBFFF800040007FFFBFFF900050006FFFAFFF900050006FFFAFFF90005",
		INIT_4F=>X"0007FFFCFFF800030007FFFCFFF800030007FFFBFFF800040007FFFBFFF80004",
		INIT_50=>X"0008FFFDFFF700020008FFFDFFF700020008FFFDFFF700020008FFFCFFF70003",
		INIT_51=>X"0008FFFFFFF700000008FFFFFFF700010008FFFEFFF700010008FFFEFFF70001",
		INIT_52=>X"00080001FFF7FFFF00080000FFF7FFFF00080000FFF7FFFF0008FFFFFFF70000",
		INIT_53=>X"00080002FFF7FFFD00080002FFF7FFFE00080001FFF7FFFE00080001FFF7FFFE",
		INIT_54=>X"00080004FFF7FFFC00080003FFF7FFFC00080003FFF7FFFC00080002FFF7FFFD",
		INIT_55=>X"00070005FFF8FFFA00070005FFF8FFFB00070004FFF8FFFB00080004FFF7FFFB",
		INIT_56=>X"00060006FFF9FFF900060006FFF9FFF900070006FFF8FFFA00070005FFF8FFFA",
		INIT_57=>X"00050007FFFAFFF800050007FFFAFFF800050007FFF9FFF800060007FFF9FFF9",
		INIT_58=>X"00030008FFFBFFF700040008FFFBFFF700040008FFFBFFF700050008FFFAFFF7",
		INIT_59=>X"00020009FFFDFFF600020009FFFCFFF600030009FFFCFFF600030009FFFCFFF7",
		INIT_5A=>X"0000000AFFFFFFF50001000AFFFEFFF600010009FFFEFFF600020009FFFDFFF6",
		INIT_5B=>X"FFFE000A0000FFF5FFFF000A0000FFF5FFFF000AFFFFFFF50000000AFFFFFFF5",
		INIT_5C=>X"FFFD000A0002FFF5FFFD000A0002FFF5FFFE000A0001FFF5FFFE000A0001FFF5",
		INIT_5D=>X"FFFB00090004FFF6FFFB00090003FFF6FFFC000A0003FFF5FFFC000A0003FFF5",
		INIT_5E=>X"FFF900090006FFF6FFFA00090005FFF6FFFA00090005FFF6FFFA00090004FFF6",
		INIT_5F=>X"FFF800080007FFF7FFF800080007FFF7FFF800080006FFF7FFF900080006FFF7",
		INIT_60=>X"FFF600060009FFF9FFF600070008FFF8FFF700070008FFF8FFF700070008FFF8",
		INIT_61=>X"FFF50005000AFFFAFFF50005000AFFFAFFF500060009FFF9FFF600060009FFF9",
		INIT_62=>X"FFF40003000BFFFCFFF40003000BFFFBFFF40004000BFFFBFFF40004000AFFFB",
		INIT_63=>X"FFF30001000CFFFEFFF30001000CFFFDFFF30002000CFFFDFFF30002000BFFFC",
		INIT_64=>X"FFF3FFFF000C0000FFF3FFFF000CFFFFFFF30000000CFFFFFFF30000000CFFFE",
		INIT_65=>X"FFF2FFFC000D0002FFF2FFFD000D0002FFF2FFFE000D0001FFF2FFFE000C0001",
		INIT_66=>X"FFF3FFFA000C0005FFF3FFFB000C0004FFF3FFFB000C0003FFF3FFFC000D0003",
		INIT_67=>X"FFF4FFF8000C0007FFF3FFF8000C0006FFF3FFF9000C0006FFF3FFF9000C0005",
		INIT_68=>X"FFF5FFF5000A0009FFF4FFF6000B0009FFF4FFF6000B0008FFF4FFF7000B0008",
		INIT_69=>X"FFF6FFF30009000CFFF6FFF40009000BFFF5FFF4000A000BFFF5FFF5000A000A",
		INIT_6A=>X"FFF8FFF10007000EFFF8FFF20008000DFFF7FFF20008000DFFF7FFF30009000C",
		INIT_6B=>X"FFFBFFEF0005000FFFFAFFF00005000FFFF9FFF00006000FFFF9FFF10007000E",
		INIT_6C=>X"FFFDFFEE00020011FFFDFFEE00030011FFFCFFEF00030010FFFBFFEF00040010",
		INIT_6D=>X"0000FFEDFFFF00120000FFED00000012FFFFFFED00010012FFFEFFEE00010011",
		INIT_6E=>X"0004FFECFFFC00130003FFECFFFC00130002FFEDFFFD00120001FFEDFFFE0012",
		INIT_6F=>X"0008FFECFFF800130007FFECFFF900130006FFECFFFA00130005FFECFFFB0013",
		INIT_70=>X"000BFFEDFFF40012000AFFECFFF500130009FFECFFF600130008FFECFFF70013",
		INIT_71=>X"000FFFEEFFF00011000EFFEDFFF10012000DFFEDFFF20012000CFFEDFFF30012",
		INIT_72=>X"0014FFF0FFEC00100013FFEFFFED00100012FFEFFFEE00110010FFEEFFEF0011",
		INIT_73=>X"0018FFF2FFE8000D0017FFF2FFE9000E0016FFF1FFEA000E0015FFF0FFEB000F",
		INIT_74=>X"001CFFF6FFE4000A001BFFF5FFE5000B001AFFF4FFE6000B0019FFF3FFE7000C",
		INIT_75=>X"0020FFFAFFDF0005001FFFF9FFE00006001EFFF8FFE10008001DFFF7FFE30009",
		INIT_76=>X"00240000FFDB00000023FFFEFFDC00010022FFFDFFDD00030021FFFCFFDE0004",
		INIT_77=>X"00280007FFD8FFF900270005FFD9FFFB00260003FFDAFFFD00250002FFDBFFFE",
		INIT_78=>X"002B0010FFD4FFF0002A000DFFD5FFF30029000BFFD6FFF500290009FFD7FFF7",
		INIT_79=>X"002E001BFFD1FFE6002E0018FFD2FFE9002D0015FFD3FFEB002C0012FFD3FFEE",
		INIT_7A=>X"00310029FFCEFFD800300025FFCFFFDC00300021FFD0FFDF002F001EFFD0FFE3",
		INIT_7B=>X"0033003DFFCCFFC500330037FFCDFFCA00320032FFCDFFCF0032002DFFCEFFD4",
		INIT_7C=>X"0035005CFFCAFFA800350052FFCBFFB10034004AFFCBFFB800340043FFCBFFBF",
		INIT_7D=>X"00360094FFC9FF7500360082FFC9FF8500360073FFC9FF9300350066FFCAFF9E",
		INIT_7E=>X"0037012DFFC8FEF3003700F2FFC8FF24003700C9FFC8FF46003700ABFFC8FF60",
		INIT_7F=>X"2038145EFFC8F93600370411FFC8FD1900370240FFC8FE290037018DFFC8FEA8",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_13,
		DOPADOP=>dopadop_13,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_14: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0",
		INITP_01=>X"3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C30F0F0F0F0",
		INITP_02=>X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F3C3C3C3C3C3C3C3C3C",
		INITP_03=>X"C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3CF0F0F0F0F0F0F0F0F0F0F0F0F0F",
		INITP_04=>X"F0F0F0F0F0F0F0F0F0F0F0F0F0F3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3",
		INITP_05=>X"3C3C3C3C3C3C3C3C3C30F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0",
		INITP_06=>X"0F0F0F0F0C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C",
		INITP_07=>X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F",
		INITP_08=>X"C30C33CF3CC30CF3CF30C33CF3CC30C33CF30C30CF3CC30C33CF3CC30CF3CF30",
		INITP_09=>X"F3CC30C33CF30C30CF3CC30C33CF3CC30CF3CF30C33CF3CC30C33CF30C30CF3C",
		INITP_0A=>X"33CF3CC30CF3CF30C33CF3CC30C33CF30C30CF3CC30C33CF3CC30CF3CF30C33C",
		INITP_0B=>X"30C33CF30C30CF3CC30C33CF3CC30CF3CF30C33CF3CC30C33CF30C30CF3CC30C",
		INITP_0C=>X"3CC30CF3CF30C30CF3CC30C33CF30C30CF3CF30C33CF3CC30CF3CF30C30CF3CC",
		INITP_0D=>X"3CF30C30CF3CF30C33CF3CC30CF3CF30C30CF3CC30C33CF30C30CF3CF30C33CF",
		INITP_0E=>X"0CF3CF30C30CF3CC30C33CF30C30CF3CF30C33CF3CC30CF3CF30C30CF3CC30C3",
		INITP_0F=>X"0C30CF3CF30C33CF3CC30CF3CF30C30CF3CC30C33CF30C30CF3CF30C33CF3CC3",
		INIT_00=>X"FFF8FFFE00070001FFF8FFFF00070000FFF8FFFF00070000FFF8FFFF00070000",
		INIT_01=>X"FFF8FFFD00070002FFF8FFFD00070002FFF8FFFE00070001FFF8FFFE00070001",
		INIT_02=>X"FFF9FFFC00070003FFF8FFFC00070003FFF8FFFC00070003FFF8FFFD00070002",
		INIT_03=>X"FFF9FFFA00060004FFF9FFFB00060004FFF9FFFB00060004FFF9FFFB00060004",
		INIT_04=>X"FFFAFFF900050005FFFAFFFA00050005FFFAFFFA00050005FFFAFFFA00060005",
		INIT_05=>X"FFFBFFF900040006FFFBFFF900040006FFFBFFF900040006FFFAFFF900050006",
		INIT_06=>X"FFFDFFF800030007FFFCFFF800030007FFFCFFF800030007FFFCFFF800040006",
		INIT_07=>X"FFFEFFF800010007FFFEFFF800020007FFFDFFF800020007FFFDFFF800020007",
		INIT_08=>X"FFFFFFF700000008FFFFFFF700000008FFFFFFF700010008FFFEFFF700010008",
		INIT_09=>X"0001FFF7FFFE00080000FFF7FFFF00080000FFF7FFFF00080000FFF700000008",
		INIT_0A=>X"0002FFF8FFFD00070002FFF8FFFD00080001FFF7FFFE00080001FFF7FFFE0008",
		INIT_0B=>X"0003FFF8FFFC00070003FFF8FFFC00070003FFF8FFFC00070002FFF8FFFD0007",
		INIT_0C=>X"0005FFF9FFFA00060004FFF9FFFB00060004FFF8FFFB00070004FFF8FFFB0007",
		INIT_0D=>X"0006FFFAFFF900050006FFF9FFFA00060005FFF9FFFA00060005FFF9FFFA0006",
		INIT_0E=>X"0007FFFBFFF800040007FFFBFFF900050006FFFAFFF900050006FFFAFFF90005",
		INIT_0F=>X"0007FFFCFFF800030007FFFCFFF800030007FFFBFFF800040007FFFBFFF80004",
		INIT_10=>X"0008FFFDFFF700020008FFFDFFF700020008FFFDFFF700020008FFFCFFF70003",
		INIT_11=>X"0008FFFFFFF700000008FFFFFFF700010008FFFEFFF700010008FFFEFFF70001",
		INIT_12=>X"00080001FFF7FFFF00080000FFF7FFFF00080000FFF7FFFF0008FFFFFFF70000",
		INIT_13=>X"00080002FFF7FFFD00080002FFF7FFFE00080001FFF7FFFE00080001FFF7FFFE",
		INIT_14=>X"00080004FFF7FFFC00080003FFF7FFFC00080003FFF7FFFC00080002FFF7FFFD",
		INIT_15=>X"00070005FFF8FFFA00070005FFF8FFFB00070004FFF8FFFB00080004FFF7FFFB",
		INIT_16=>X"00060006FFF9FFF900060006FFF9FFF900070006FFF8FFFA00070005FFF8FFFA",
		INIT_17=>X"00050007FFFAFFF800050007FFFAFFF800050007FFF9FFF800060007FFF9FFF9",
		INIT_18=>X"00030008FFFBFFF700040008FFFBFFF700040008FFFBFFF700050008FFFAFFF7",
		INIT_19=>X"00020009FFFDFFF600020009FFFCFFF600030009FFFCFFF600030009FFFCFFF7",
		INIT_1A=>X"0000000AFFFFFFF50001000AFFFEFFF600010009FFFEFFF600020009FFFDFFF6",
		INIT_1B=>X"FFFE000A0000FFF5FFFF000A0000FFF5FFFF000AFFFFFFF50000000AFFFFFFF5",
		INIT_1C=>X"FFFD000A0002FFF5FFFD000A0002FFF5FFFE000A0001FFF5FFFE000A0001FFF5",
		INIT_1D=>X"FFFB00090004FFF6FFFB00090003FFF6FFFC000A0003FFF5FFFC000A0003FFF5",
		INIT_1E=>X"FFF900090006FFF6FFFA00090005FFF6FFFA00090005FFF6FFFA00090004FFF6",
		INIT_1F=>X"FFF800080007FFF7FFF800080007FFF7FFF800080006FFF7FFF900080006FFF7",
		INIT_20=>X"FFF600060009FFF9FFF600070008FFF8FFF700070008FFF8FFF700070008FFF8",
		INIT_21=>X"FFF50005000AFFFAFFF50005000AFFFAFFF500060009FFF9FFF600060009FFF9",
		INIT_22=>X"FFF40003000BFFFCFFF40003000BFFFBFFF40004000BFFFBFFF40004000AFFFB",
		INIT_23=>X"FFF30001000CFFFEFFF30001000CFFFDFFF30002000CFFFDFFF30002000BFFFC",
		INIT_24=>X"FFF3FFFF000C0000FFF3FFFF000CFFFFFFF30000000CFFFFFFF30000000CFFFE",
		INIT_25=>X"FFF2FFFC000D0002FFF2FFFD000D0002FFF2FFFE000D0001FFF2FFFE000C0001",
		INIT_26=>X"FFF3FFFA000C0005FFF3FFFB000C0004FFF3FFFB000C0003FFF3FFFC000D0003",
		INIT_27=>X"FFF4FFF8000C0007FFF3FFF8000C0006FFF3FFF9000C0006FFF3FFF9000C0005",
		INIT_28=>X"FFF5FFF5000A0009FFF4FFF6000B0009FFF4FFF6000B0008FFF4FFF7000B0008",
		INIT_29=>X"FFF6FFF30009000CFFF6FFF40009000BFFF5FFF4000A000BFFF5FFF5000A000A",
		INIT_2A=>X"FFF8FFF10007000EFFF8FFF20008000DFFF7FFF20008000DFFF7FFF30009000C",
		INIT_2B=>X"FFFBFFEF0005000FFFFAFFF00005000FFFF9FFF00006000FFFF9FFF10007000E",
		INIT_2C=>X"FFFDFFEE00020011FFFDFFEE00030011FFFCFFEF00030010FFFBFFEF00040010",
		INIT_2D=>X"0000FFEDFFFF00120000FFED00000012FFFFFFED00010012FFFEFFEE00010011",
		INIT_2E=>X"0004FFECFFFC00130003FFECFFFC00130002FFEDFFFD00120001FFEDFFFE0012",
		INIT_2F=>X"0008FFECFFF800130007FFECFFF900130006FFECFFFA00130005FFECFFFB0013",
		INIT_30=>X"000BFFEDFFF40012000AFFECFFF500130009FFECFFF600130008FFECFFF70013",
		INIT_31=>X"000FFFEEFFF00011000EFFEDFFF10012000DFFEDFFF20012000CFFEDFFF30012",
		INIT_32=>X"0014FFF0FFEC00100013FFEFFFED00100012FFEFFFEE00110010FFEEFFEF0011",
		INIT_33=>X"0018FFF2FFE8000D0017FFF2FFE9000E0016FFF1FFEA000E0015FFF0FFEB000F",
		INIT_34=>X"001CFFF6FFE4000A001BFFF5FFE5000B001AFFF4FFE6000B0019FFF3FFE7000C",
		INIT_35=>X"0020FFFAFFDF0005001FFFF9FFE00006001EFFF8FFE10008001DFFF7FFE30009",
		INIT_36=>X"00240000FFDB00000023FFFEFFDC00010022FFFDFFDD00030021FFFCFFDE0004",
		INIT_37=>X"00280007FFD8FFF900270005FFD9FFFB00260003FFDAFFFD00250002FFDBFFFE",
		INIT_38=>X"002B0010FFD4FFF0002A000DFFD5FFF30029000BFFD6FFF500290009FFD7FFF7",
		INIT_39=>X"002E001BFFD1FFE6002E0018FFD2FFE9002D0015FFD3FFEB002C0012FFD3FFEE",
		INIT_3A=>X"00310029FFCEFFD800300025FFCFFFDC00300021FFD0FFDF002F001EFFD0FFE3",
		INIT_3B=>X"0033003DFFCCFFC500330037FFCDFFCA00320032FFCDFFCF0032002DFFCEFFD4",
		INIT_3C=>X"0035005CFFCAFFA800350052FFCBFFB10034004AFFCBFFB800340043FFCBFFBF",
		INIT_3D=>X"00360094FFC9FF7500360082FFC9FF8500360073FFC9FF9300350066FFCAFF9E",
		INIT_3E=>X"0037012DFFC8FEF3003700F2FFC8FF24003700C9FFC8FF46003700ABFFC8FF60",
		INIT_3F=>X"2038145EFFC8F93600370411FFC8FD1900370240FFC8FE290037018DFFC8FEA8",
		INIT_40=>X"00050001FFF80007FFFEFFFA0007FFFCFFFC0007FFF9FFFF0006FFF800020004",
		INIT_41=>X"0001FFF80007FFFEFFFA0007FFFBFFFD0007FFF9FFFF0006FFF800020004FFF8",
		INIT_42=>X"FFF90007FFFDFFFB0008FFFBFFFD0007FFF900000006FFF800030003FFF80005",
		INIT_43=>X"0007FFFDFFFB0008FFFAFFFE0007FFF800010005FFF800030003FFF800060000",
		INIT_44=>X"FFFCFFFC0007FFFAFFFE0007FFF800010005FFF700040002FFF800060000FFF9",
		INIT_45=>X"FFFC0007FFF9FFFF0006FFF800020004FFF700040002FFF80006FFFFFFF90007",
		INIT_46=>X"0007FFF9FFFF0006FFF800020004FFF700050001FFF80007FFFEFFFA0007FFFC",
		INIT_47=>X"FFF900000006FFF800030004FFF700050001FFF80007FFFEFFFA0008FFFBFFFD",
		INIT_48=>X"00010005FFF700030003FFF700060000FFF90007FFFDFFFA0008FFFBFFFD0007",
		INIT_49=>X"0005FFF700040003FFF800060000FFF90007FFFDFFFB0008FFFAFFFE0007FFF8",
		INIT_4A=>X"FFF700040002FFF80006FFFFFFF90008FFFCFFFB0008FFFAFFFE0007FFF80001",
		INIT_4B=>X"00050001FFF80007FFFFFFF90008FFFCFFFC0008FFF9FFFF0007FFF800020005",
		INIT_4C=>X"0001FFF80007FFFEFFFA0008FFFBFFFC0008FFF9FFFF0006FFF800020004FFF7",
		INIT_4D=>X"FFF80007FFFDFFFA0008FFFBFFFD0008FFF900000006FFF700030004FFF70005",
		INIT_4E=>X"0008FFFDFFFB0008FFFAFFFD0007FFF800000006FFF700030003FFF700060000",
		INIT_4F=>X"FFFCFFFB0008FFFAFFFE0007FFF800010005FFF700040003FFF700060000FFF8",
		INIT_50=>X"FFFC0008FFF9FFFF0007FFF700020005FFF700040002FFF70007FFFFFFF90008",
		INIT_51=>X"0008FFF9FFFF0007FFF700020005FFF700050002FFF70007FFFFFFF90008FFFC",
		INIT_52=>X"FFF800000006FFF700030004FFF700060001FFF80007FFFEFFF90008FFFBFFFC",
		INIT_53=>X"00000006FFF700030004FFF700060001FFF80008FFFDFFFA0008FFFAFFFD0008",
		INIT_54=>X"0006FFF600040003FFF700070000FFF80008FFFDFFFA0009FFFAFFFD0008FFF8",
		INIT_55=>X"FFF600050003FFF70007FFFFFFF80008FFFCFFFB0009FFF9FFFE0008FFF70001",
		INIT_56=>X"00050002FFF70008FFFFFFF90009FFFBFFFB0009FFF9FFFE0008FFF700020005",
		INIT_57=>X"0001FFF70008FFFEFFF90009FFFBFFFC0009FFF8FFFF0007FFF700020005FFF6",
		INIT_58=>X"FFF70008FFFDFFF90009FFFAFFFC0009FFF800000007FFF600030005FFF60006",
		INIT_59=>X"0009FFFDFFFA0009FFF9FFFD0009FFF700000007FFF600040004FFF600070001",
		INIT_5A=>X"FFFCFFFA000AFFF9FFFD0009FFF700010007FFF600040004FFF600070000FFF7",
		INIT_5B=>X"FFFB000AFFF8FFFE0008FFF600020006FFF500050003FFF60008FFFFFFF70009",
		INIT_5C=>X"000AFFF7FFFF0008FFF600030006FFF500060002FFF60008FFFFFFF8000AFFFB",
		INIT_5D=>X"FFF700000008FFF500030005FFF500070002FFF60009FFFEFFF8000AFFFAFFFB",
		INIT_5E=>X"00000008FFF500040005FFF500070001FFF60009FFFDFFF8000AFFFAFFFC000A",
		INIT_5F=>X"0008FFF400050004FFF500080000FFF6000AFFFCFFF9000BFFF9FFFC000AFFF6",
		INIT_60=>X"FFF400060004FFF400090000FFF6000BFFFCFFF9000BFFF8FFFD000AFFF60001",
		INIT_61=>X"00070003FFF40009FFFFFFF7000BFFFBFFFA000BFFF7FFFE000AFFF500020007",
		INIT_62=>X"0002FFF4000AFFFEFFF7000CFFFAFFFA000BFFF6FFFF000AFFF400030007FFF4",
		INIT_63=>X"FFF4000BFFFDFFF7000CFFF9FFFB000BFFF6FFFF0009FFF400040006FFF30007",
		INIT_64=>X"000CFFFCFFF8000CFFF8FFFC000CFFF500000009FFF300050006FFF300080001",
		INIT_65=>X"FFFBFFF8000DFFF7FFFD000CFFF400010009FFF200060005FFF300090001FFF4",
		INIT_66=>X"FFF9000DFFF6FFFD000CFFF300020009FFF200070004FFF2000A0000FFF5000C",
		INIT_67=>X"000EFFF5FFFE000CFFF200030008FFF100080004FFF2000BFFFFFFF5000DFFFA",
		INIT_68=>X"FFF4FFFF000CFFF100040008FFF100090003FFF2000CFFFEFFF5000EFFF9FFF9",
		INIT_69=>X"0000000BFFF000060007FFF0000A0002FFF2000DFFFDFFF5000FFFF8FFFA000E",
		INIT_6A=>X"000BFFF000070007FFF0000B0001FFF2000EFFFBFFF6000FFFF6FFFB000EFFF3",
		INIT_6B=>X"FFEF00080006FFEF000D0000FFF2000FFFFAFFF60010FFF5FFFC000FFFF10001",
		INIT_6C=>X"000A0005FFEF000EFFFFFFF20010FFF9FFF70011FFF4FFFD000FFFF00003000B",
		INIT_6D=>X"0004FFEE0010FFFDFFF20012FFF7FFF70011FFF2FFFE000FFFEF0004000BFFEE",
		INIT_6E=>X"FFEE0011FFFCFFF20013FFF6FFF80012FFF1FFFF000FFFED0006000AFFED000B",
		INIT_6F=>X"0013FFFAFFF20014FFF4FFF90013FFEF0000000FFFEC0007000AFFEC000D0003",
		INIT_70=>X"FFF9FFF30016FFF2FFFA0014FFED0002000FFFEA00090009FFEB000F0002FFED",
		INIT_71=>X"FFF30017FFF0FFFB0014FFEB0004000FFFE9000B0008FFEA00110000FFED0015",
		INIT_72=>X"0019FFEDFFFD0015FFE80006000FFFE7000D0007FFE80013FFFFFFED0017FFF6",
		INIT_73=>X"FFEAFFFE0016FFE60008000FFFE500100006FFE70016FFFDFFEC0019FFF4FFF4",
		INIT_74=>X"00000017FFE3000A000FFFE200130005FFE60019FFFBFFEC001BFFF1FFF5001A",
		INIT_75=>X"0018FFDF000E000EFFE000170003FFE4001CFFF8FFEC001EFFEEFFF6001CFFE7",
		INIT_76=>X"FFDB0012000EFFDD001B0001FFE20020FFF5FFEB0022FFEBFFF7001FFFE30003",
		INIT_77=>X"0016000DFFD90020FFFFFFE00025FFF1FFEB0026FFE6FFF80021FFDE00050019",
		INIT_78=>X"000CFFD40027FFFCFFDE002BFFECFFEB002BFFE0FFFA0025FFD90009001AFFD6",
		INIT_79=>X"FFCE002FFFF7FFDB0033FFE6FFEB0031FFD9FFFD0029FFD1000E001CFFD0001C",
		INIT_7A=>X"003BFFF1FFD6003EFFDDFFEB003AFFCF0000002EFFC80014001EFFC70025000A",
		INIT_7B=>X"FFE8FFD0004FFFD0FFEB0046FFC000050036FFB9001E0020FFBC00300008FFC6",
		INIT_7C=>X"FFC5006AFFBBFFEA005BFFA9000E0042FFA3002C0024FFA900420005FFB9004D",
		INIT_7D=>X"00A1FF8FFFEA0082FF7B001E0059FF7A0047002BFF880061FFFFFFA3006DFFD8",
		INIT_7E=>X"FF09FFEA00F3FEFE004A0094FF120088003CFF3C00A9FFF1FF7300AFFFB7FFAF",
		INIT_7F=>X"2D18104EF639026002C0FBEF0239009DFDAF01FCFFB5FEB101AEFF3FFF650153",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_14,
		DOPADOP=>dopadop_14,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
	mem_15: RAMB36E1 generic map (
		READ_WIDTH_A=>18,
		INITP_00=>X"C30C33CF3CC30CF3CF30C33CF3CC30C33CF30C30CF3CC30C33CF3CC30CF3CF30",
		INITP_01=>X"F3CC30C33CF30C30CF3CC30C33CF3CC30CF3CF30C33CF3CC30C33CF30C30CF3C",
		INITP_02=>X"33CF3CC30CF3CF30C33CF3CC30C33CF30C30CF3CC30C33CF3CC30CF3CF30C33C",
		INITP_03=>X"30C33CF30C30CF3CC30C33CF3CC30CF3CF30C33CF3CC30C33CF30C30CF3CC30C",
		INITP_04=>X"3CC30CF3CF30C30CF3CC30C33CF30C30CF3CF30C33CF3CC30CF3CF30C30CF3CC",
		INITP_05=>X"3CF30C30CF3CF30C33CF3CC30CF3CF30C30CF3CC30C33CF30C30CF3CF30C33CF",
		INITP_06=>X"0CF3CF30C30CF3CC30C33CF30C30CF3CF30C33CF3CC30CF3CF30C30CF3CC30C3",
		INITP_07=>X"0C30CF3CF30C33CF3CC30CF3CF30C30CF3CC30C33CF30C30CF3CF30C33CF3CC3",
		INITP_08=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_09=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000",
		INITP_0A=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0B=>X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0C=>X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_0D=>X"FFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000",
		INITP_0E=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INITP_0F=>X"3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_00=>X"00050001FFF80007FFFEFFFA0007FFFCFFFC0007FFF9FFFF0006FFF800020004",
		INIT_01=>X"0001FFF80007FFFEFFFA0007FFFBFFFD0007FFF9FFFF0006FFF800020004FFF8",
		INIT_02=>X"FFF90007FFFDFFFB0008FFFBFFFD0007FFF900000006FFF800030003FFF80005",
		INIT_03=>X"0007FFFDFFFB0008FFFAFFFE0007FFF800010005FFF800030003FFF800060000",
		INIT_04=>X"FFFCFFFC0007FFFAFFFE0007FFF800010005FFF700040002FFF800060000FFF9",
		INIT_05=>X"FFFC0007FFF9FFFF0006FFF800020004FFF700040002FFF80006FFFFFFF90007",
		INIT_06=>X"0007FFF9FFFF0006FFF800020004FFF700050001FFF80007FFFEFFFA0007FFFC",
		INIT_07=>X"FFF900000006FFF800030004FFF700050001FFF80007FFFEFFFA0008FFFBFFFD",
		INIT_08=>X"00010005FFF700030003FFF700060000FFF90007FFFDFFFA0008FFFBFFFD0007",
		INIT_09=>X"0005FFF700040003FFF800060000FFF90007FFFDFFFB0008FFFAFFFE0007FFF8",
		INIT_0A=>X"FFF700040002FFF80006FFFFFFF90008FFFCFFFB0008FFFAFFFE0007FFF80001",
		INIT_0B=>X"00050001FFF80007FFFFFFF90008FFFCFFFC0008FFF9FFFF0007FFF800020005",
		INIT_0C=>X"0001FFF80007FFFEFFFA0008FFFBFFFC0008FFF9FFFF0006FFF800020004FFF7",
		INIT_0D=>X"FFF80007FFFDFFFA0008FFFBFFFD0008FFF900000006FFF700030004FFF70005",
		INIT_0E=>X"0008FFFDFFFB0008FFFAFFFD0007FFF800000006FFF700030003FFF700060000",
		INIT_0F=>X"FFFCFFFB0008FFFAFFFE0007FFF800010005FFF700040003FFF700060000FFF8",
		INIT_10=>X"FFFC0008FFF9FFFF0007FFF700020005FFF700040002FFF70007FFFFFFF90008",
		INIT_11=>X"0008FFF9FFFF0007FFF700020005FFF700050002FFF70007FFFFFFF90008FFFC",
		INIT_12=>X"FFF800000006FFF700030004FFF700060001FFF80007FFFEFFF90008FFFBFFFC",
		INIT_13=>X"00000006FFF700030004FFF700060001FFF80008FFFDFFFA0008FFFAFFFD0008",
		INIT_14=>X"0006FFF600040003FFF700070000FFF80008FFFDFFFA0009FFFAFFFD0008FFF8",
		INIT_15=>X"FFF600050003FFF70007FFFFFFF80008FFFCFFFB0009FFF9FFFE0008FFF70001",
		INIT_16=>X"00050002FFF70008FFFFFFF90009FFFBFFFB0009FFF9FFFE0008FFF700020005",
		INIT_17=>X"0001FFF70008FFFEFFF90009FFFBFFFC0009FFF8FFFF0007FFF700020005FFF6",
		INIT_18=>X"FFF70008FFFDFFF90009FFFAFFFC0009FFF800000007FFF600030005FFF60006",
		INIT_19=>X"0009FFFDFFFA0009FFF9FFFD0009FFF700000007FFF600040004FFF600070001",
		INIT_1A=>X"FFFCFFFA000AFFF9FFFD0009FFF700010007FFF600040004FFF600070000FFF7",
		INIT_1B=>X"FFFB000AFFF8FFFE0008FFF600020006FFF500050003FFF60008FFFFFFF70009",
		INIT_1C=>X"000AFFF7FFFF0008FFF600030006FFF500060002FFF60008FFFFFFF8000AFFFB",
		INIT_1D=>X"FFF700000008FFF500030005FFF500070002FFF60009FFFEFFF8000AFFFAFFFB",
		INIT_1E=>X"00000008FFF500040005FFF500070001FFF60009FFFDFFF8000AFFFAFFFC000A",
		INIT_1F=>X"0008FFF400050004FFF500080000FFF6000AFFFCFFF9000BFFF9FFFC000AFFF6",
		INIT_20=>X"FFF400060004FFF400090000FFF6000BFFFCFFF9000BFFF8FFFD000AFFF60001",
		INIT_21=>X"00070003FFF40009FFFFFFF7000BFFFBFFFA000BFFF7FFFE000AFFF500020007",
		INIT_22=>X"0002FFF4000AFFFEFFF7000CFFFAFFFA000BFFF6FFFF000AFFF400030007FFF4",
		INIT_23=>X"FFF4000BFFFDFFF7000CFFF9FFFB000BFFF6FFFF0009FFF400040006FFF30007",
		INIT_24=>X"000CFFFCFFF8000CFFF8FFFC000CFFF500000009FFF300050006FFF300080001",
		INIT_25=>X"FFFBFFF8000DFFF7FFFD000CFFF400010009FFF200060005FFF300090001FFF4",
		INIT_26=>X"FFF9000DFFF6FFFD000CFFF300020009FFF200070004FFF2000A0000FFF5000C",
		INIT_27=>X"000EFFF5FFFE000CFFF200030008FFF100080004FFF2000BFFFFFFF5000DFFFA",
		INIT_28=>X"FFF4FFFF000CFFF100040008FFF100090003FFF2000CFFFEFFF5000EFFF9FFF9",
		INIT_29=>X"0000000BFFF000060007FFF0000A0002FFF2000DFFFDFFF5000FFFF8FFFA000E",
		INIT_2A=>X"000BFFF000070007FFF0000B0001FFF2000EFFFBFFF6000FFFF6FFFB000EFFF3",
		INIT_2B=>X"FFEF00080006FFEF000D0000FFF2000FFFFAFFF60010FFF5FFFC000FFFF10001",
		INIT_2C=>X"000A0005FFEF000EFFFFFFF20010FFF9FFF70011FFF4FFFD000FFFF00003000B",
		INIT_2D=>X"0004FFEE0010FFFDFFF20012FFF7FFF70011FFF2FFFE000FFFEF0004000BFFEE",
		INIT_2E=>X"FFEE0011FFFCFFF20013FFF6FFF80012FFF1FFFF000FFFED0006000AFFED000B",
		INIT_2F=>X"0013FFFAFFF20014FFF4FFF90013FFEF0000000FFFEC0007000AFFEC000D0003",
		INIT_30=>X"FFF9FFF30016FFF2FFFA0014FFED0002000FFFEA00090009FFEB000F0002FFED",
		INIT_31=>X"FFF30017FFF0FFFB0014FFEB0004000FFFE9000B0008FFEA00110000FFED0015",
		INIT_32=>X"0019FFEDFFFD0015FFE80006000FFFE7000D0007FFE80013FFFFFFED0017FFF6",
		INIT_33=>X"FFEAFFFE0016FFE60008000FFFE500100006FFE70016FFFDFFEC0019FFF4FFF4",
		INIT_34=>X"00000017FFE3000A000FFFE200130005FFE60019FFFBFFEC001BFFF1FFF5001A",
		INIT_35=>X"0018FFDF000E000EFFE000170003FFE4001CFFF8FFEC001EFFEEFFF6001CFFE7",
		INIT_36=>X"FFDB0012000EFFDD001B0001FFE20020FFF5FFEB0022FFEBFFF7001FFFE30003",
		INIT_37=>X"0016000DFFD90020FFFFFFE00025FFF1FFEB0026FFE6FFF80021FFDE00050019",
		INIT_38=>X"000CFFD40027FFFCFFDE002BFFECFFEB002BFFE0FFFA0025FFD90009001AFFD6",
		INIT_39=>X"FFCE002FFFF7FFDB0033FFE6FFEB0031FFD9FFFD0029FFD1000E001CFFD0001C",
		INIT_3A=>X"003BFFF1FFD6003EFFDDFFEB003AFFCF0000002EFFC80014001EFFC70025000A",
		INIT_3B=>X"FFE8FFD0004FFFD0FFEB0046FFC000050036FFB9001E0020FFBC00300008FFC6",
		INIT_3C=>X"FFC5006AFFBBFFEA005BFFA9000E0042FFA3002C0024FFA900420005FFB9004D",
		INIT_3D=>X"00A1FF8FFFEA0082FF7B001E0059FF7A0047002BFF880061FFFFFFA3006DFFD8",
		INIT_3E=>X"FF09FFEA00F3FEFE004A0094FF120088003CFF3C00A9FFF1FF7300AFFFB7FFAF",
		INIT_3F=>X"2D18104EF639026002C0FBEF0239009DFDAF01FCFFB5FEB101AEFF3FFF650153",
		INIT_40=>X"0007000700070007000700070007000700070007000700070007000700070007",
		INIT_41=>X"0007000700070007000700070007000700070007000700070007000700070007",
		INIT_42=>X"0006000700070007000700070007000700070007000700070007000700070007",
		INIT_43=>X"0006000600060006000600060006000600060006000600060006000600060006",
		INIT_44=>X"0005000500050005000500050005000500050005000500050005000600060006",
		INIT_45=>X"0004000400040004000400040004000400040004000400040005000500050005",
		INIT_46=>X"0002000300030003000300030003000300030003000300030003000300040004",
		INIT_47=>X"0001000100010001000100020002000200020002000200020002000200020002",
		INIT_48=>X"0000000000000000000000000000000000000000000100010001000100010001",
		INIT_49=>X"FFFEFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000",
		INIT_4A=>X"FFFDFFFDFFFDFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFE",
		INIT_4B=>X"FFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFD",
		INIT_4C=>X"FFFAFFFAFFFAFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFB",
		INIT_4D=>X"FFF9FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFA",
		INIT_4E=>X"FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_4F=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_50=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_51=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_52=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_53=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_54=>X"FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7FFF7",
		INIT_55=>X"FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF7FFF7FFF7FFF7FFF7",
		INIT_56=>X"FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8",
		INIT_57=>X"FFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFFAFFF9FFF9FFF9FFF9FFF9FFF9FFF9",
		INIT_58=>X"FFFCFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFBFFFAFFFAFFFAFFFA",
		INIT_59=>X"FFFDFFFDFFFDFFFDFFFDFFFDFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFC",
		INIT_5A=>X"FFFFFFFFFFFFFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFEFFFDFFFDFFFDFFFD",
		INIT_5B=>X"0001000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_5C=>X"0002000200020002000200020002000200010001000100010001000100010001",
		INIT_5D=>X"0004000400040004000400040003000300030003000300030003000300030002",
		INIT_5E=>X"0006000600060006000500050005000500050005000500050005000400040004",
		INIT_5F=>X"0008000700070007000700070007000700070007000600060006000600060006",
		INIT_60=>X"0009000900090009000900090008000800080008000800080008000800080008",
		INIT_61=>X"000A000A000A000A000A000A000A000A000A000A000900090009000900090009",
		INIT_62=>X"000B000B000B000B000B000B000B000B000B000B000B000B000B000A000A000A",
		INIT_63=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000B000B000B",
		INIT_64=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C",
		INIT_65=>X"000D000D000D000D000D000D000D000D000D000D000D000D000D000D000C000C",
		INIT_66=>X"000C000C000C000C000C000C000C000C000C000C000C000C000C000C000D000D",
		INIT_67=>X"000B000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C",
		INIT_68=>X"000A000A000A000B000B000B000B000B000B000B000B000B000B000B000B000B",
		INIT_69=>X"0009000900090009000900090009000A000A000A000A000A000A000A000A000A",
		INIT_6A=>X"0007000700070007000700070008000800080008000800080008000800090009",
		INIT_6B=>X"0004000500050005000500050005000600060006000600060006000600070007",
		INIT_6C=>X"0002000200020002000200030003000300030003000300040004000400040004",
		INIT_6D=>X"FFFFFFFFFFFFFFFFFFFF00000000000000000000000100010001000100010001",
		INIT_6E=>X"FFFBFFFBFFFCFFFCFFFCFFFCFFFCFFFDFFFDFFFDFFFDFFFEFFFEFFFEFFFEFFFE",
		INIT_6F=>X"FFF8FFF8FFF8FFF8FFF8FFF9FFF9FFF9FFF9FFFAFFFAFFFAFFFAFFFBFFFBFFFB",
		INIT_70=>X"FFF4FFF4FFF4FFF4FFF5FFF5FFF5FFF5FFF6FFF6FFF6FFF6FFF7FFF7FFF7FFF7",
		INIT_71=>X"FFF0FFF0FFF0FFF0FFF1FFF1FFF1FFF1FFF2FFF2FFF2FFF2FFF3FFF3FFF3FFF3",
		INIT_72=>X"FFEBFFECFFECFFECFFECFFEDFFEDFFEDFFEDFFEEFFEEFFEEFFEFFFEFFFEFFFEF",
		INIT_73=>X"FFE7FFE7FFE8FFE8FFE8FFE9FFE9FFE9FFE9FFEAFFEAFFEAFFEAFFEBFFEBFFEB",
		INIT_74=>X"FFE3FFE3FFE4FFE4FFE4FFE4FFE5FFE5FFE5FFE5FFE6FFE6FFE6FFE6FFE7FFE7",
		INIT_75=>X"FFDFFFDFFFDFFFE0FFE0FFE0FFE0FFE1FFE1FFE1FFE1FFE2FFE2FFE2FFE3FFE3",
		INIT_76=>X"FFDBFFDBFFDBFFDCFFDCFFDCFFDCFFDDFFDDFFDDFFDDFFDEFFDEFFDEFFDEFFDF",
		INIT_77=>X"FFD7FFD8FFD8FFD8FFD8FFD8FFD9FFD9FFD9FFD9FFDAFFDAFFDAFFDAFFDBFFDB",
		INIT_78=>X"FFD4FFD4FFD4FFD4FFD5FFD5FFD5FFD5FFD6FFD6FFD6FFD6FFD6FFD7FFD7FFD7",
		INIT_79=>X"FFD1FFD1FFD1FFD1FFD1FFD2FFD2FFD2FFD2FFD2FFD3FFD3FFD3FFD3FFD3FFD4",
		INIT_7A=>X"FFCEFFCEFFCEFFCEFFCFFFCFFFCFFFCFFFCFFFCFFFD0FFD0FFD0FFD0FFD0FFD1",
		INIT_7B=>X"FFCCFFCCFFCCFFCCFFCCFFCCFFCDFFCDFFCDFFCDFFCDFFCDFFCDFFCEFFCEFFCE",
		INIT_7C=>X"FFCAFFCAFFCAFFCAFFCAFFCAFFCBFFCBFFCBFFCBFFCBFFCBFFCBFFCBFFCBFFCC",
		INIT_7D=>X"FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFC9FFCAFFCAFFCAFFCA",
		INIT_7E=>X"FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC9",
		INIT_7F=>X"3FC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8FFC8",
		SIM_DEVICE=>"7SERIES"
	)port map(
		CASCADEOUTA=>open,
		CASCADEOUTB=>open,
		DBITERR=>open,
		ECCPARITY=>open,
		RDADDRECC=>open,
		SBITERR=>open,
		DOADO=>doado_15,
		DOPADOP=>dopadop_15,
		DOBDO=>open,
		DOPBDOP=>open,
		CASCADEINA=>'0',
		CASCADEINB=>'0',
		INJECTDBITERR=>'0',
		INJECTSBITERR=>'0',
		ADDRARDADDR=>addrardaddr,
		CLKARDCLK=>clk,
		ENARDEN=>'1',
		REGCEAREGCE=>'1',
		RSTRAMARSTRAM=>'0',
		RSTREGARSTREG=>'0',
		WEA=>b"0000",
		DIADI=>(others=>'0'),
		DIPADIP=>(others=>'0'),
		ADDRBWRADDR=>(others=>'0'),
		CLKBWRCLK=>'0',
		ENBWREN=>'0',
		REGCEB=>'0',
		RSTRAMB=>'0',
		RSTREGB=>'0',
		WEBWE=>(others=>'0'),
		DIBDI=>(others=>'0'),
		DIPBDIP=>(others=>'0')
	);
end arch;
